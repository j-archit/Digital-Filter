`timescale 1ns / 1ps

module testbench;

    // Parameters and Inputs
    parameter htp = 10;   // Half time Period of Clock
    reg clk, reset;
    reg signed [31:0] x;
    wire signed [31:0] y;

    // Instantiate the Unit Under Test (DUT)
    iir_N #(.N(2)) DUT(
      .clk(clk),
      .rst(reset),
      .x(x),
      .y(y)
    );

    // Generate clock with 100ns period
    initial clk = 0;
    always #htp clk = ~clk;
    
    always @(posedge(clk)) begin
      $display("%.0f,%.0f", x, y);
    end
    

    initial begin
        x = 32'd0;
        reset = 1;
        clk = 0;
        clk = 1;
        #10;
        reset = 0;
        #20;

        x =               25; #(2*htp); // Sample(1)
        x =               10; #(2*htp); // Sample(1)
        x =               25; #(2*htp); // Sample(1)
        x =               10; #(2*htp); // Sample(1)
        x =               67; #(2*htp); // Sample(1)
        x =              -56; #(2*htp); // Sample(2)
        x =               19; #(2*htp); // Sample(3)
        x =               28; #(2*htp); // Sample(4)
        x =              160; #(2*htp); // Sample(5)
        x =               39; #(2*htp); // Sample(6)
        x =              142; #(2*htp); // Sample(7)
        x =              151; #(2*htp); // Sample(8)
        x =              117; #(2*htp); // Sample(9)
        x =              294; #(2*htp); // Sample(10)
        x =              199; #(2*htp); // Sample(11)
        x =              363; #(2*htp); // Sample(12)
        x =              100; #(2*htp); // Sample(13)
        x =              525; #(2*htp); // Sample(14)
        x =               78; #(2*htp); // Sample(15)
        x =              195; #(2*htp); // Sample(16)
        x =              -19; #(2*htp); // Sample(17)
        x =              147; #(2*htp); // Sample(18)
        x =              515; #(2*htp); // Sample(19)
        x =              373; #(2*htp); // Sample(20)
        x =              110; #(2*htp); // Sample(21)
        x =              389; #(2*htp); // Sample(22)
        x =              161; #(2*htp); // Sample(23)
        x =              -98; #(2*htp); // Sample(24)
        x =              198; #(2*htp); // Sample(25)
        x =              673; #(2*htp); // Sample(26)
        x =              338; #(2*htp); // Sample(27)
        x =              -79; #(2*htp); // Sample(28)
        x =              424; #(2*htp); // Sample(29)
        x =              653; #(2*htp); // Sample(30)
        x =              269; #(2*htp); // Sample(31)
        x =              241; #(2*htp); // Sample(32)
        x =              374; #(2*htp); // Sample(33)
        x =               92; #(2*htp); // Sample(34)
        x =              296; #(2*htp); // Sample(35)
        x =              707; #(2*htp); // Sample(36)
        x =               46; #(2*htp); // Sample(37)
        x =              212; #(2*htp); // Sample(38)
        x =              262; #(2*htp); // Sample(39)
        x =              251; #(2*htp); // Sample(40)
        x =              315; #(2*htp); // Sample(41)
        x =               94; #(2*htp); // Sample(42)
        x =              -26; #(2*htp); // Sample(43)
        x =               84; #(2*htp); // Sample(44)
        x =             -286; #(2*htp); // Sample(45)
        x =               18; #(2*htp); // Sample(46)
        x =              459; #(2*htp); // Sample(47)
        x =              -86; #(2*htp); // Sample(48)
        x =               70; #(2*htp); // Sample(49)
        x =               77; #(2*htp); // Sample(50)
        x =               38; #(2*htp); // Sample(51)
        x =              -44; #(2*htp); // Sample(52)
        x =             -200; #(2*htp); // Sample(53)
        x =              -27; #(2*htp); // Sample(54)
        x =              -67; #(2*htp); // Sample(55)
        x =             -100; #(2*htp); // Sample(56)
        x =              -33; #(2*htp); // Sample(57)
        x =             -199; #(2*htp); // Sample(58)
        x =             -407; #(2*htp); // Sample(59)
        x =             -343; #(2*htp); // Sample(60)
        x =              -78; #(2*htp); // Sample(61)
        x =              -28; #(2*htp); // Sample(62)
        x =             -358; #(2*htp); // Sample(63)
        x =             -503; #(2*htp); // Sample(64)
        x =             -454; #(2*htp); // Sample(65)
        x =              -75; #(2*htp); // Sample(66)
        x =             -101; #(2*htp); // Sample(67)
        x =             -133; #(2*htp); // Sample(68)
        x =             -103; #(2*htp); // Sample(69)
        x =             -299; #(2*htp); // Sample(70)
        x =             -267; #(2*htp); // Sample(71)
        x =             -161; #(2*htp); // Sample(72)
        x =             -123; #(2*htp); // Sample(73)
        x =              191; #(2*htp); // Sample(74)
        x =             -482; #(2*htp); // Sample(75)
        x =             -272; #(2*htp); // Sample(76)
        x =             -206; #(2*htp); // Sample(77)
        x =             -506; #(2*htp); // Sample(78)
        x =             -562; #(2*htp); // Sample(79)
        x =             -238; #(2*htp); // Sample(80)
        x =             -396; #(2*htp); // Sample(81)
        x =             -249; #(2*htp); // Sample(82)
        x =             -421; #(2*htp); // Sample(83)
        x =             -245; #(2*htp); // Sample(84)
        x =             -193; #(2*htp); // Sample(85)
        x =             -624; #(2*htp); // Sample(86)
        x =              -37; #(2*htp); // Sample(87)
        x =             -554; #(2*htp); // Sample(88)
        x =             -101; #(2*htp); // Sample(89)
        x =             -129; #(2*htp); // Sample(90)
        x =              -70; #(2*htp); // Sample(91)
        x =              197; #(2*htp); // Sample(92)
        x =             -374; #(2*htp); // Sample(93)
        x =             -191; #(2*htp); // Sample(94)
        x =             -186; #(2*htp); // Sample(95)
        x =              278; #(2*htp); // Sample(96)
        x =              253; #(2*htp); // Sample(97)
        x =              156; #(2*htp); // Sample(98)
        x =             -260; #(2*htp); // Sample(99)
        x =              -30; #(2*htp); // Sample(100)
        x =              179; #(2*htp); // Sample(101)
        x =              164; #(2*htp); // Sample(102)
        x =              -10; #(2*htp); // Sample(103)
        x =              423; #(2*htp); // Sample(104)
        x =               39; #(2*htp); // Sample(105)
        x =              241; #(2*htp); // Sample(106)
        x =              568; #(2*htp); // Sample(107)
        x =              532; #(2*htp); // Sample(108)
        x =              174; #(2*htp); // Sample(109)
        x =              371; #(2*htp); // Sample(110)
        x =              562; #(2*htp); // Sample(111)
        x =               66; #(2*htp); // Sample(112)
        x =              445; #(2*htp); // Sample(113)
        x =              628; #(2*htp); // Sample(114)
        x =              471; #(2*htp); // Sample(115)
        x =              522; #(2*htp); // Sample(116)
        x =              290; #(2*htp); // Sample(117)
        x =               47; #(2*htp); // Sample(118)
        x =              157; #(2*htp); // Sample(119)
        x =              597; #(2*htp); // Sample(120)
        x =              314; #(2*htp); // Sample(121)
        x =              458; #(2*htp); // Sample(122)
        x =              102; #(2*htp); // Sample(123)
        x =              -47; #(2*htp); // Sample(124)
        x =             -105; #(2*htp); // Sample(125)
        x =              338; #(2*htp); // Sample(126)
        x =             -133; #(2*htp); // Sample(127)
        x =              543; #(2*htp); // Sample(128)
        x =              479; #(2*htp); // Sample(129)
        x =              307; #(2*htp); // Sample(130)
        x =              435; #(2*htp); // Sample(131)
        x =              206; #(2*htp); // Sample(132)
        x =             -133; #(2*htp); // Sample(133)
        x =              174; #(2*htp); // Sample(134)
        x =               55; #(2*htp); // Sample(135)
        x =              405; #(2*htp); // Sample(136)
        x =              216; #(2*htp); // Sample(137)
        x =              211; #(2*htp); // Sample(138)
        x =               45; #(2*htp); // Sample(139)
        x =              -72; #(2*htp); // Sample(140)
        x =              131; #(2*htp); // Sample(141)
        x =              -23; #(2*htp); // Sample(142)
        x =              301; #(2*htp); // Sample(143)
        x =              -49; #(2*htp); // Sample(144)
        x =             -150; #(2*htp); // Sample(145)
        x =              -61; #(2*htp); // Sample(146)
        x =              165; #(2*htp); // Sample(147)
        x =             -166; #(2*htp); // Sample(148)
        x =              -96; #(2*htp); // Sample(149)
        x =             -374; #(2*htp); // Sample(150)
        x =              -92; #(2*htp); // Sample(151)
        x =             -205; #(2*htp); // Sample(152)
        x =             -234; #(2*htp); // Sample(153)
        x =             -140; #(2*htp); // Sample(154)
        x =             -178; #(2*htp); // Sample(155)
        x =             -198; #(2*htp); // Sample(156)
        x =              354; #(2*htp); // Sample(157)
        x =              -29; #(2*htp); // Sample(158)
        x =               80; #(2*htp); // Sample(159)
        x =               65; #(2*htp); // Sample(160)
        x =             -314; #(2*htp); // Sample(161)
        x =             -361; #(2*htp); // Sample(162)
        x =             -591; #(2*htp); // Sample(163)
        x =             -467; #(2*htp); // Sample(164)
        x =             -344; #(2*htp); // Sample(165)
        x =             -311; #(2*htp); // Sample(166)
        x =             -236; #(2*htp); // Sample(167)
        x =             -270; #(2*htp); // Sample(168)
        x =             -525; #(2*htp); // Sample(169)
        x =             -361; #(2*htp); // Sample(170)
        x =               30; #(2*htp); // Sample(171)
        x =             -351; #(2*htp); // Sample(172)
        x =             -464; #(2*htp); // Sample(173)
        x =             -332; #(2*htp); // Sample(174)
        x =             -214; #(2*htp); // Sample(175)
        x =             -342; #(2*htp); // Sample(176)
        x =             -341; #(2*htp); // Sample(177)
        x =             -314; #(2*htp); // Sample(178)
        x =              -13; #(2*htp); // Sample(179)
        x =              -67; #(2*htp); // Sample(180)
        x =             -354; #(2*htp); // Sample(181)
        x =             -339; #(2*htp); // Sample(182)
        x =             -512; #(2*htp); // Sample(183)
        x =               46; #(2*htp); // Sample(184)
        x =             -170; #(2*htp); // Sample(185)
        x =             -179; #(2*htp); // Sample(186)
        x =              -81; #(2*htp); // Sample(187)
        x =             -342; #(2*htp); // Sample(188)
        x =             -252; #(2*htp); // Sample(189)
        x =              -24; #(2*htp); // Sample(190)
        x =             -100; #(2*htp); // Sample(191)
        x =             -409; #(2*htp); // Sample(192)
        x =             -146; #(2*htp); // Sample(193)
        x =               70; #(2*htp); // Sample(194)
        x =              242; #(2*htp); // Sample(195)
        x =               76; #(2*htp); // Sample(196)
        x =              105; #(2*htp); // Sample(197)
        x =                5; #(2*htp); // Sample(198)
        x =              155; #(2*htp); // Sample(199)
        x =              236; #(2*htp); // Sample(200)
        x =              -21; #(2*htp); // Sample(201)
        x =              366; #(2*htp); // Sample(202)
        x =             -132; #(2*htp); // Sample(203)
        x =              189; #(2*htp); // Sample(204)
        x =              168; #(2*htp); // Sample(205)
        x =              538; #(2*htp); // Sample(206)
        x =              179; #(2*htp); // Sample(207)
        x =              861; #(2*htp); // Sample(208)
        x =              208; #(2*htp); // Sample(209)
        x =              133; #(2*htp); // Sample(210)
        x =              718; #(2*htp); // Sample(211)
        x =              280; #(2*htp); // Sample(212)
        x =              241; #(2*htp); // Sample(213)
        x =              322; #(2*htp); // Sample(214)
        x =              107; #(2*htp); // Sample(215)
        x =               22; #(2*htp); // Sample(216)
        x =              178; #(2*htp); // Sample(217)
        x =              312; #(2*htp); // Sample(218)
        x =              514; #(2*htp); // Sample(219)
        x =              524; #(2*htp); // Sample(220)
        x =              381; #(2*htp); // Sample(221)
        x =              511; #(2*htp); // Sample(222)
        x =              775; #(2*htp); // Sample(223)
        x =              393; #(2*htp); // Sample(224)
        x =              443; #(2*htp); // Sample(225)
        x =              192; #(2*htp); // Sample(226)
        x =              466; #(2*htp); // Sample(227)
        x =               12; #(2*htp); // Sample(228)
        x =              149; #(2*htp); // Sample(229)
        x =               35; #(2*htp); // Sample(230)
        x =               77; #(2*htp); // Sample(231)
        x =              545; #(2*htp); // Sample(232)
        x =              111; #(2*htp); // Sample(233)
        x =               52; #(2*htp); // Sample(234)
        x =              311; #(2*htp); // Sample(235)
        x =               36; #(2*htp); // Sample(236)
        x =              139; #(2*htp); // Sample(237)
        x =              164; #(2*htp); // Sample(238)
        x =             -126; #(2*htp); // Sample(239)
        x =              -47; #(2*htp); // Sample(240)
        x =              365; #(2*htp); // Sample(241)
        x =                6; #(2*htp); // Sample(242)
        x =              133; #(2*htp); // Sample(243)
        x =              184; #(2*htp); // Sample(244)
        x =               32; #(2*htp); // Sample(245)
        x =              -72; #(2*htp); // Sample(246)
        x =              129; #(2*htp); // Sample(247)
        x =             -372; #(2*htp); // Sample(248)
        x =               80; #(2*htp); // Sample(249)
        x =             -567; #(2*htp); // Sample(250)
        x =             -423; #(2*htp); // Sample(251)
        x =             -279; #(2*htp); // Sample(252)
        x =             -228; #(2*htp); // Sample(253)
        x =             -536; #(2*htp); // Sample(254)
        x =              -90; #(2*htp); // Sample(255)
        x =             -264; #(2*htp); // Sample(256)
        x =             -469; #(2*htp); // Sample(257)
        x =             -496; #(2*htp); // Sample(258)
        x =             -460; #(2*htp); // Sample(259)
        x =             -443; #(2*htp); // Sample(260)
        x =             -314; #(2*htp); // Sample(261)
        x =             -304; #(2*htp); // Sample(262)
        x =             -408; #(2*htp); // Sample(263)
        x =             -315; #(2*htp); // Sample(264)
        x =             -423; #(2*htp); // Sample(265)
        x =             -265; #(2*htp); // Sample(266)
        x =               -2; #(2*htp); // Sample(267)
        x =             -130; #(2*htp); // Sample(268)
        x =             -368; #(2*htp); // Sample(269)
        x =             -256; #(2*htp); // Sample(270)
        x =             -307; #(2*htp); // Sample(271)
        x =             -350; #(2*htp); // Sample(272)
        x =             -320; #(2*htp); // Sample(273)
        x =              -38; #(2*htp); // Sample(274)
        x =             -342; #(2*htp); // Sample(275)
        x =             -190; #(2*htp); // Sample(276)
        x =              -95; #(2*htp); // Sample(277)
        x =             -395; #(2*htp); // Sample(278)
        x =             -470; #(2*htp); // Sample(279)
        x =              -21; #(2*htp); // Sample(280)
        x =              -77; #(2*htp); // Sample(281)
        x =             -235; #(2*htp); // Sample(282)
        x =              100; #(2*htp); // Sample(283)
        x =              -36; #(2*htp); // Sample(284)
        x =             -155; #(2*htp); // Sample(285)
        x =             -143; #(2*htp); // Sample(286)
        x =             -134; #(2*htp); // Sample(287)
        x =             -228; #(2*htp); // Sample(288)
        x =              519; #(2*htp); // Sample(289)
        x =             -412; #(2*htp); // Sample(290)
        x =               91; #(2*htp); // Sample(291)
        x =               60; #(2*htp); // Sample(292)
        x =             -166; #(2*htp); // Sample(293)
        x =               68; #(2*htp); // Sample(294)
        x =              189; #(2*htp); // Sample(295)
        x =              328; #(2*htp); // Sample(296)
        x =              171; #(2*htp); // Sample(297)
        x =              278; #(2*htp); // Sample(298)
        x =              516; #(2*htp); // Sample(299)
        x =              177; #(2*htp); // Sample(300)
        x =              103; #(2*htp); // Sample(301)
        x =              -46; #(2*htp); // Sample(302)
        x =              399; #(2*htp); // Sample(303)
        x =              152; #(2*htp); // Sample(304)
        x =              530; #(2*htp); // Sample(305)
        x =              283; #(2*htp); // Sample(306)
        x =              251; #(2*htp); // Sample(307)
        x =              177; #(2*htp); // Sample(308)
        x =              192; #(2*htp); // Sample(309)
        x =               54; #(2*htp); // Sample(310)
        x =              411; #(2*htp); // Sample(311)
        x =              219; #(2*htp); // Sample(312)
        x =              421; #(2*htp); // Sample(313)
        x =              -22; #(2*htp); // Sample(314)
        x =              362; #(2*htp); // Sample(315)
        x =              120; #(2*htp); // Sample(316)
        x =               -7; #(2*htp); // Sample(317)
        x =              239; #(2*htp); // Sample(318)
        x =              394; #(2*htp); // Sample(319)
        x =              465; #(2*htp); // Sample(320)
        x =              494; #(2*htp); // Sample(321)
        x =              177; #(2*htp); // Sample(322)
        x =               56; #(2*htp); // Sample(323)
        x =              802; #(2*htp); // Sample(324)
        x =              108; #(2*htp); // Sample(325)
        x =               64; #(2*htp); // Sample(326)
        x =              273; #(2*htp); // Sample(327)
        x =              -37; #(2*htp); // Sample(328)
        x =               24; #(2*htp); // Sample(329)
        x =             -156; #(2*htp); // Sample(330)
        x =               77; #(2*htp); // Sample(331)
        x =             -117; #(2*htp); // Sample(332)
        x =              152; #(2*htp); // Sample(333)
        x =               95; #(2*htp); // Sample(334)
        x =              -97; #(2*htp); // Sample(335)
        x =              -53; #(2*htp); // Sample(336)
        x =             -108; #(2*htp); // Sample(337)
        x =               12; #(2*htp); // Sample(338)
        x =             -163; #(2*htp); // Sample(339)
        x =               -8; #(2*htp); // Sample(340)
        x =             -239; #(2*htp); // Sample(341)
        x =               15; #(2*htp); // Sample(342)
        x =             -146; #(2*htp); // Sample(343)
        x =             -521; #(2*htp); // Sample(344)
        x =             -114; #(2*htp); // Sample(345)
        x =               12; #(2*htp); // Sample(346)
        x =               56; #(2*htp); // Sample(347)
        x =             -155; #(2*htp); // Sample(348)
        x =               68; #(2*htp); // Sample(349)
        x =              -95; #(2*htp); // Sample(350)
        x =              160; #(2*htp); // Sample(351)
        x =             -199; #(2*htp); // Sample(352)
        x =             -169; #(2*htp); // Sample(353)
        x =             -187; #(2*htp); // Sample(354)
        x =             -172; #(2*htp); // Sample(355)
        x =             -127; #(2*htp); // Sample(356)
        x =              -89; #(2*htp); // Sample(357)
        x =             -480; #(2*htp); // Sample(358)
        x =             -542; #(2*htp); // Sample(359)
        x =              -47; #(2*htp); // Sample(360)
        x =             -117; #(2*htp); // Sample(361)
        x =             -459; #(2*htp); // Sample(362)
        x =             -306; #(2*htp); // Sample(363)
        x =               55; #(2*htp); // Sample(364)
        x =             -508; #(2*htp); // Sample(365)
        x =             -222; #(2*htp); // Sample(366)
        x =             -539; #(2*htp); // Sample(367)
        x =             -236; #(2*htp); // Sample(368)
        x =             -202; #(2*htp); // Sample(369)
        x =             -283; #(2*htp); // Sample(370)
        x =              -60; #(2*htp); // Sample(371)
        x =             -252; #(2*htp); // Sample(372)
        x =               12; #(2*htp); // Sample(373)
        x =                9; #(2*htp); // Sample(374)
        x =             -235; #(2*htp); // Sample(375)
        x =             -118; #(2*htp); // Sample(376)
        x =             -110; #(2*htp); // Sample(377)
        x =               50; #(2*htp); // Sample(378)
        x =              120; #(2*htp); // Sample(379)
        x =               54; #(2*htp); // Sample(380)
        x =              -73; #(2*htp); // Sample(381)
        x =             -227; #(2*htp); // Sample(382)
        x =             -282; #(2*htp); // Sample(383)
        x =              188; #(2*htp); // Sample(384)
        x =              377; #(2*htp); // Sample(385)
        x =               71; #(2*htp); // Sample(386)
        x =               26; #(2*htp); // Sample(387)
        x =              236; #(2*htp); // Sample(388)
        x =             -239; #(2*htp); // Sample(389)
        x =               47; #(2*htp); // Sample(390)
        x =             -262; #(2*htp); // Sample(391)
        x =              214; #(2*htp); // Sample(392)
        x =              156; #(2*htp); // Sample(393)
        x =              229; #(2*htp); // Sample(394)
        x =              102; #(2*htp); // Sample(395)
        x =             -154; #(2*htp); // Sample(396)
        x =              400; #(2*htp); // Sample(397)
        x =              103; #(2*htp); // Sample(398)
        x =              272; #(2*htp); // Sample(399)
        x =              429; #(2*htp); // Sample(400)
        x =              368; #(2*htp); // Sample(401)
        x =              113; #(2*htp); // Sample(402)
        x =              228; #(2*htp); // Sample(403)
        x =              243; #(2*htp); // Sample(404)
        x =              477; #(2*htp); // Sample(405)
        x =              537; #(2*htp); // Sample(406)
        x =               97; #(2*htp); // Sample(407)
        x =              107; #(2*htp); // Sample(408)
        x =              325; #(2*htp); // Sample(409)
        x =              299; #(2*htp); // Sample(410)
        x =              335; #(2*htp); // Sample(411)
        x =               96; #(2*htp); // Sample(412)
        x =               37; #(2*htp); // Sample(413)
        x =              269; #(2*htp); // Sample(414)
        x =              511; #(2*htp); // Sample(415)
        x =              389; #(2*htp); // Sample(416)
        x =              238; #(2*htp); // Sample(417)
        x =              177; #(2*htp); // Sample(418)
        x =               26; #(2*htp); // Sample(419)
        x =              396; #(2*htp); // Sample(420)
        x =              374; #(2*htp); // Sample(421)
        x =              167; #(2*htp); // Sample(422)
        x =              256; #(2*htp); // Sample(423)
        x =              219; #(2*htp); // Sample(424)
        x =              325; #(2*htp); // Sample(425)
        x =              443; #(2*htp); // Sample(426)
        x =             -217; #(2*htp); // Sample(427)
        x =               38; #(2*htp); // Sample(428)
        x =               63; #(2*htp); // Sample(429)
        x =             -182; #(2*htp); // Sample(430)
        x =              -16; #(2*htp); // Sample(431)
        x =              174; #(2*htp); // Sample(432)
        x =             -143; #(2*htp); // Sample(433)
        x =             -417; #(2*htp); // Sample(434)
        x =             -232; #(2*htp); // Sample(435)
        x =               -5; #(2*htp); // Sample(436)
        x =             -222; #(2*htp); // Sample(437)
        x =               83; #(2*htp); // Sample(438)
        x =             -220; #(2*htp); // Sample(439)
        x =              -89; #(2*htp); // Sample(440)
        x =             -263; #(2*htp); // Sample(441)
        x =              -48; #(2*htp); // Sample(442)
        x =             -493; #(2*htp); // Sample(443)
        x =              112; #(2*htp); // Sample(444)
        x =             -253; #(2*htp); // Sample(445)
        x =             -252; #(2*htp); // Sample(446)
        x =             -507; #(2*htp); // Sample(447)
        x =             -249; #(2*htp); // Sample(448)
        x =             -273; #(2*htp); // Sample(449)
        x =             -497; #(2*htp); // Sample(450)
        x =             -164; #(2*htp); // Sample(451)
        x =               96; #(2*htp); // Sample(452)
        x =              -65; #(2*htp); // Sample(453)
        x =             -306; #(2*htp); // Sample(454)
        x =             -192; #(2*htp); // Sample(455)
        x =             -259; #(2*htp); // Sample(456)
        x =             -221; #(2*htp); // Sample(457)
        x =             -689; #(2*htp); // Sample(458)
        x =             -468; #(2*htp); // Sample(459)
        x =             -348; #(2*htp); // Sample(460)
        x =             -170; #(2*htp); // Sample(461)
        x =             -215; #(2*htp); // Sample(462)
        x =             -296; #(2*htp); // Sample(463)
        x =             -677; #(2*htp); // Sample(464)
        x =             -529; #(2*htp); // Sample(465)
        x =                4; #(2*htp); // Sample(466)
        x =             -212; #(2*htp); // Sample(467)
        x =             -223; #(2*htp); // Sample(468)
        x =             -276; #(2*htp); // Sample(469)
        x =              351; #(2*htp); // Sample(470)
        x =             -312; #(2*htp); // Sample(471)
        x =             -194; #(2*htp); // Sample(472)
        x =              -49; #(2*htp); // Sample(473)
        x =              117; #(2*htp); // Sample(474)
        x =             -140; #(2*htp); // Sample(475)
        x =               87; #(2*htp); // Sample(476)
        x =              110; #(2*htp); // Sample(477)
        x =              -10; #(2*htp); // Sample(478)
        x =             -287; #(2*htp); // Sample(479)
        x =              132; #(2*htp); // Sample(480)
        x =               20; #(2*htp); // Sample(481)
        x =              313; #(2*htp); // Sample(482)
        x =             -119; #(2*htp); // Sample(483)
        x =               58; #(2*htp); // Sample(484)
        x =              -17; #(2*htp); // Sample(485)
        x =             -251; #(2*htp); // Sample(486)
        x =              -83; #(2*htp); // Sample(487)
        x =             -236; #(2*htp); // Sample(488)
        x =              469; #(2*htp); // Sample(489)
        x =              213; #(2*htp); // Sample(490)
        x =              296; #(2*htp); // Sample(491)
        x =              237; #(2*htp); // Sample(492)
        x =              423; #(2*htp); // Sample(493)
        x =              512; #(2*htp); // Sample(494)
        x =              162; #(2*htp); // Sample(495)
        x =               67; #(2*htp); // Sample(496)
        x =              469; #(2*htp); // Sample(497)
        x =              693; #(2*htp); // Sample(498)
        x =              236; #(2*htp); // Sample(499)
        x =              141; #(2*htp); // Sample(500)
        x =                0; #(2*htp); // Sample(1)
        x =              183; #(2*htp); // Sample(2)
        x =              290; #(2*htp); // Sample(3)
        x =              277; #(2*htp); // Sample(4)
        x =              150; #(2*htp); // Sample(5)
        x =              -39; #(2*htp); // Sample(6)
        x =             -212; #(2*htp); // Sample(7)
        x =             -297; #(2*htp); // Sample(8)
        x =             -260; #(2*htp); // Sample(9)
        x =             -115; #(2*htp); // Sample(10)
        x =               78; #(2*htp); // Sample(11)
        x =              238; #(2*htp); // Sample(12)
        x =              300; #(2*htp); // Sample(13)
        x =              238; #(2*htp); // Sample(14)
        x =               78; #(2*htp); // Sample(15)
        x =             -115; #(2*htp); // Sample(16)
        x =             -260; #(2*htp); // Sample(17)
        x =             -297; #(2*htp); // Sample(18)
        x =             -212; #(2*htp); // Sample(19)
        x =              -39; #(2*htp); // Sample(20)
        x =              150; #(2*htp); // Sample(21)
        x =              277; #(2*htp); // Sample(22)
        x =              290; #(2*htp); // Sample(23)
        x =              183; #(2*htp); // Sample(24)
        x =                0; #(2*htp); // Sample(25)
        x =             -183; #(2*htp); // Sample(26)
        x =             -290; #(2*htp); // Sample(27)
        x =             -277; #(2*htp); // Sample(28)
        x =             -150; #(2*htp); // Sample(29)
        x =               39; #(2*htp); // Sample(30)
        x =              212; #(2*htp); // Sample(31)
        x =              297; #(2*htp); // Sample(32)
        x =              260; #(2*htp); // Sample(33)
        x =              115; #(2*htp); // Sample(34)
        x =              -78; #(2*htp); // Sample(35)
        x =             -238; #(2*htp); // Sample(36)
        x =             -300; #(2*htp); // Sample(37)
        x =             -238; #(2*htp); // Sample(38)
        x =              -78; #(2*htp); // Sample(39)
        x =              115; #(2*htp); // Sample(40)
        x =              260; #(2*htp); // Sample(41)
        x =              297; #(2*htp); // Sample(42)
        x =              212; #(2*htp); // Sample(43)
        x =               39; #(2*htp); // Sample(44)
        x =             -150; #(2*htp); // Sample(45)
        x =             -277; #(2*htp); // Sample(46)
        x =             -290; #(2*htp); // Sample(47)
        x =             -183; #(2*htp); // Sample(48)
        x =               -0; #(2*htp); // Sample(49)
        x =              183; #(2*htp); // Sample(50)
        x =              290; #(2*htp); // Sample(51)
        x =              277; #(2*htp); // Sample(52)

/*
        x =              150; #(2*htp); // Sample(53)
        x =              -39; #(2*htp); // Sample(54)
        x =             -212; #(2*htp); // Sample(55)
        x =             -297; #(2*htp); // Sample(56)
        x =             -260; #(2*htp); // Sample(57)
        x =             -115; #(2*htp); // Sample(58)
        x =               78; #(2*htp); // Sample(59)
        x =              238; #(2*htp); // Sample(60)
        x =              300; #(2*htp); // Sample(61)
        x =              238; #(2*htp); // Sample(62)
        x =               78; #(2*htp); // Sample(63)
        x =             -115; #(2*htp); // Sample(64)
        x =             -260; #(2*htp); // Sample(65)
        x =             -297; #(2*htp); // Sample(66)
        x =             -212; #(2*htp); // Sample(67)
        x =              -39; #(2*htp); // Sample(68)
        x =              150; #(2*htp); // Sample(69)
        x =              277; #(2*htp); // Sample(70)
        x =              290; #(2*htp); // Sample(71)
        x =              183; #(2*htp); // Sample(72)
        x =               -0; #(2*htp); // Sample(73)
        x =             -183; #(2*htp); // Sample(74)
        x =             -290; #(2*htp); // Sample(75)
        x =             -277; #(2*htp); // Sample(76)
        x =             -150; #(2*htp); // Sample(77)
        x =               39; #(2*htp); // Sample(78)
        x =              212; #(2*htp); // Sample(79)
        x =              297; #(2*htp); // Sample(80)
        x =              260; #(2*htp); // Sample(81)
        x =              115; #(2*htp); // Sample(82)
        x =              -78; #(2*htp); // Sample(83)
        x =             -238; #(2*htp); // Sample(84)
        x =             -300; #(2*htp); // Sample(85)
        x =             -238; #(2*htp); // Sample(86)
        x =              -78; #(2*htp); // Sample(87)
        x =              115; #(2*htp); // Sample(88)
        x =              260; #(2*htp); // Sample(89)
        x =              297; #(2*htp); // Sample(90)
        x =              212; #(2*htp); // Sample(91)
        x =               39; #(2*htp); // Sample(92)
        x =             -150; #(2*htp); // Sample(93)
        x =             -277; #(2*htp); // Sample(94)
        x =             -290; #(2*htp); // Sample(95)
        x =             -183; #(2*htp); // Sample(96)
        x =               -0; #(2*htp); // Sample(97)
        x =              183; #(2*htp); // Sample(98)
        x =              290; #(2*htp); // Sample(99)
        x =              277; #(2*htp); // Sample(100)
        x =              150; #(2*htp); // Sample(101)
        x =              -39; #(2*htp); // Sample(102)
        x =             -212; #(2*htp); // Sample(103)
        x =             -297; #(2*htp); // Sample(104)
        x =             -260; #(2*htp); // Sample(105)
        x =             -115; #(2*htp); // Sample(106)
        x =               78; #(2*htp); // Sample(107)
        x =              238; #(2*htp); // Sample(108)
        x =              300; #(2*htp); // Sample(109)
        x =              238; #(2*htp); // Sample(110)
        x =               78; #(2*htp); // Sample(111)
        x =             -115; #(2*htp); // Sample(112)
        x =             -260; #(2*htp); // Sample(113)
        x =             -297; #(2*htp); // Sample(114)
        x =             -212; #(2*htp); // Sample(115)
        x =              -39; #(2*htp); // Sample(116)
        x =              150; #(2*htp); // Sample(117)
        x =              277; #(2*htp); // Sample(118)
        x =              290; #(2*htp); // Sample(119)
        x =              183; #(2*htp); // Sample(120)
        x =               -0; #(2*htp); // Sample(121)
        x =             -183; #(2*htp); // Sample(122)
        x =             -290; #(2*htp); // Sample(123)
        x =             -277; #(2*htp); // Sample(124)
        x =             -150; #(2*htp); // Sample(125)
        x =               39; #(2*htp); // Sample(126)
        x =              212; #(2*htp); // Sample(127)
        x =              297; #(2*htp); // Sample(128)
        x =              260; #(2*htp); // Sample(129)
        x =              115; #(2*htp); // Sample(130)
        x =              -78; #(2*htp); // Sample(131)
        x =             -238; #(2*htp); // Sample(132)
        x =             -300; #(2*htp); // Sample(133)
        x =             -238; #(2*htp); // Sample(134)
        x =              -78; #(2*htp); // Sample(135)
        x =              115; #(2*htp); // Sample(136)
        x =              260; #(2*htp); // Sample(137)
        x =              297; #(2*htp); // Sample(138)
        x =              212; #(2*htp); // Sample(139)
        x =               39; #(2*htp); // Sample(140)
        x =             -150; #(2*htp); // Sample(141)
        x =             -277; #(2*htp); // Sample(142)
        x =             -290; #(2*htp); // Sample(143)
        x =             -183; #(2*htp); // Sample(144)
        x =                0; #(2*htp); // Sample(145)
        x =              183; #(2*htp); // Sample(146)
        x =              290; #(2*htp); // Sample(147)
        x =              277; #(2*htp); // Sample(148)
        x =              150; #(2*htp); // Sample(149)
        x =              -39; #(2*htp); // Sample(150)
        x =             -212; #(2*htp); // Sample(151)
        x =             -297; #(2*htp); // Sample(152)
        x =             -260; #(2*htp); // Sample(153)
        x =             -115; #(2*htp); // Sample(154)
        x =               78; #(2*htp); // Sample(155)
        x =              238; #(2*htp); // Sample(156)
        x =              300; #(2*htp); // Sample(157)
        x =              238; #(2*htp); // Sample(158)
        x =               78; #(2*htp); // Sample(159)
        x =             -115; #(2*htp); // Sample(160)
        x =             -260; #(2*htp); // Sample(161)
        x =             -297; #(2*htp); // Sample(162)
        x =             -212; #(2*htp); // Sample(163)
        x =              -39; #(2*htp); // Sample(164)
        x =              150; #(2*htp); // Sample(165)
        x =              277; #(2*htp); // Sample(166)
        x =              290; #(2*htp); // Sample(167)
        x =              183; #(2*htp); // Sample(168)
        x =               -0; #(2*htp); // Sample(169)
        x =             -183; #(2*htp); // Sample(170)
        x =             -290; #(2*htp); // Sample(171)
        x =             -277; #(2*htp); // Sample(172)
        x =             -150; #(2*htp); // Sample(173)
        x =               39; #(2*htp); // Sample(174)
        x =              212; #(2*htp); // Sample(175)
        x =              297; #(2*htp); // Sample(176)
        x =              260; #(2*htp); // Sample(177)
        x =              115; #(2*htp); // Sample(178)
        x =              -78; #(2*htp); // Sample(179)
        x =             -238; #(2*htp); // Sample(180)
        x =             -300; #(2*htp); // Sample(181)
        x =             -238; #(2*htp); // Sample(182)
        x =              -78; #(2*htp); // Sample(183)
        x =              115; #(2*htp); // Sample(184)
        x =              260; #(2*htp); // Sample(185)
        x =              297; #(2*htp); // Sample(186)
        x =              212; #(2*htp); // Sample(187)
        x =               39; #(2*htp); // Sample(188)
        x =             -150; #(2*htp); // Sample(189)
        x =             -277; #(2*htp); // Sample(190)
        x =             -290; #(2*htp); // Sample(191)
        x =             -183; #(2*htp); // Sample(192)
        x =               -0; #(2*htp); // Sample(193)
        x =              183; #(2*htp); // Sample(194)
        x =              290; #(2*htp); // Sample(195)
        x =              277; #(2*htp); // Sample(196)
        x =              150; #(2*htp); // Sample(197)
        x =              -39; #(2*htp); // Sample(198)
        x =             -212; #(2*htp); // Sample(199)
        x =             -297; #(2*htp); // Sample(200)
        x =             -260; #(2*htp); // Sample(201)
        x =             -115; #(2*htp); // Sample(202)
        x =               78; #(2*htp); // Sample(203)
        x =              238; #(2*htp); // Sample(204)
        x =              300; #(2*htp); // Sample(205)
        x =              238; #(2*htp); // Sample(206)
        x =               78; #(2*htp); // Sample(207)
        x =             -115; #(2*htp); // Sample(208)
        x =             -260; #(2*htp); // Sample(209)
        x =             -297; #(2*htp); // Sample(210)
        x =             -212; #(2*htp); // Sample(211)
        x =              -39; #(2*htp); // Sample(212)
        x =              150; #(2*htp); // Sample(213)
        x =              277; #(2*htp); // Sample(214)
        x =              290; #(2*htp); // Sample(215)
        x =              183; #(2*htp); // Sample(216)
        x =                0; #(2*htp); // Sample(217)
        x =             -183; #(2*htp); // Sample(218)
        x =             -290; #(2*htp); // Sample(219)
        x =             -277; #(2*htp); // Sample(220)
        x =             -150; #(2*htp); // Sample(221)
        x =               39; #(2*htp); // Sample(222)
        x =              212; #(2*htp); // Sample(223)
        x =              297; #(2*htp); // Sample(224)
        x =              260; #(2*htp); // Sample(225)
        x =              115; #(2*htp); // Sample(226)
        x =              -78; #(2*htp); // Sample(227)
        x =             -238; #(2*htp); // Sample(228)
        x =             -300; #(2*htp); // Sample(229)
        x =             -238; #(2*htp); // Sample(230)
        x =              -78; #(2*htp); // Sample(231)
        x =              115; #(2*htp); // Sample(232)
        x =              260; #(2*htp); // Sample(233)
        x =              297; #(2*htp); // Sample(234)
        x =              212; #(2*htp); // Sample(235)
        x =               39; #(2*htp); // Sample(236)
        x =             -150; #(2*htp); // Sample(237)
        x =             -277; #(2*htp); // Sample(238)
        x =             -290; #(2*htp); // Sample(239)
        x =             -183; #(2*htp); // Sample(240)
        x =                0; #(2*htp); // Sample(241)
        x =              183; #(2*htp); // Sample(242)
        x =              290; #(2*htp); // Sample(243)
        x =              277; #(2*htp); // Sample(244)
        x =              150; #(2*htp); // Sample(245)
        x =              -39; #(2*htp); // Sample(246)
        x =             -212; #(2*htp); // Sample(247)
        x =             -297; #(2*htp); // Sample(248)
        x =             -260; #(2*htp); // Sample(249)
        x =             -115; #(2*htp); // Sample(250)
        x =               78; #(2*htp); // Sample(251)
        x =              238; #(2*htp); // Sample(252)
        x =              300; #(2*htp); // Sample(253)
        x =              238; #(2*htp); // Sample(254)
        x =               78; #(2*htp); // Sample(255)
        x =             -115; #(2*htp); // Sample(256)
        x =             -260; #(2*htp); // Sample(257)
        x =             -297; #(2*htp); // Sample(258)
        x =             -212; #(2*htp); // Sample(259)
        x =              -39; #(2*htp); // Sample(260)
        x =              150; #(2*htp); // Sample(261)
        x =              277; #(2*htp); // Sample(262)
        x =              290; #(2*htp); // Sample(263)
        x =              183; #(2*htp); // Sample(264)
        x =               -0; #(2*htp); // Sample(265)
        x =             -183; #(2*htp); // Sample(266)
        x =             -290; #(2*htp); // Sample(267)
        x =             -277; #(2*htp); // Sample(268)
        x =             -150; #(2*htp); // Sample(269)
        x =               39; #(2*htp); // Sample(270)
        x =              212; #(2*htp); // Sample(271)
        x =              297; #(2*htp); // Sample(272)
        x =              260; #(2*htp); // Sample(273)
        x =              115; #(2*htp); // Sample(274)
        x =              -78; #(2*htp); // Sample(275)
        x =             -238; #(2*htp); // Sample(276)
        x =             -300; #(2*htp); // Sample(277)
        x =             -238; #(2*htp); // Sample(278)
        x =              -78; #(2*htp); // Sample(279)
        x =              115; #(2*htp); // Sample(280)
        x =              260; #(2*htp); // Sample(281)
        x =              297; #(2*htp); // Sample(282)
        x =              212; #(2*htp); // Sample(283)
        x =               39; #(2*htp); // Sample(284)
        x =             -150; #(2*htp); // Sample(285)
        x =             -277; #(2*htp); // Sample(286)
        x =             -290; #(2*htp); // Sample(287)
        x =             -183; #(2*htp); // Sample(288)
        x =                0; #(2*htp); // Sample(289)
        x =              183; #(2*htp); // Sample(290)
        x =              290; #(2*htp); // Sample(291)
        x =              277; #(2*htp); // Sample(292)
        x =              150; #(2*htp); // Sample(293)
        x =              -39; #(2*htp); // Sample(294)
        x =             -212; #(2*htp); // Sample(295)
        x =             -297; #(2*htp); // Sample(296)
        x =             -260; #(2*htp); // Sample(297)
        x =             -115; #(2*htp); // Sample(298)
        x =               78; #(2*htp); // Sample(299)
        x =              238; #(2*htp); // Sample(300)
        x =              300; #(2*htp); // Sample(301)
        x =              238; #(2*htp); // Sample(302)
        x =               78; #(2*htp); // Sample(303)
        x =             -115; #(2*htp); // Sample(304)
        x =             -260; #(2*htp); // Sample(305)
        x =             -297; #(2*htp); // Sample(306)
        x =             -212; #(2*htp); // Sample(307)
        x =              -39; #(2*htp); // Sample(308)
        x =              150; #(2*htp); // Sample(309)
        x =              277; #(2*htp); // Sample(310)
        x =              290; #(2*htp); // Sample(311)
        x =              183; #(2*htp); // Sample(312)
        x =               -0; #(2*htp); // Sample(313)
        x =             -183; #(2*htp); // Sample(314)
        x =             -290; #(2*htp); // Sample(315)
        x =             -277; #(2*htp); // Sample(316)
        x =             -150; #(2*htp); // Sample(317)
        x =               39; #(2*htp); // Sample(318)
        x =              212; #(2*htp); // Sample(319)
        x =              297; #(2*htp); // Sample(320)
        x =              260; #(2*htp); // Sample(321)
        x =              115; #(2*htp); // Sample(322)
        x =              -78; #(2*htp); // Sample(323)
        x =             -238; #(2*htp); // Sample(324)
        x =             -300; #(2*htp); // Sample(325)
        x =             -238; #(2*htp); // Sample(326)
        x =              -78; #(2*htp); // Sample(327)
        x =              115; #(2*htp); // Sample(328)
        x =              260; #(2*htp); // Sample(329)
        x =              297; #(2*htp); // Sample(330)
        x =              212; #(2*htp); // Sample(331)
        x =               39; #(2*htp); // Sample(332)
        x =             -150; #(2*htp); // Sample(333)
        x =             -277; #(2*htp); // Sample(334)
        x =             -290; #(2*htp); // Sample(335)
        x =             -183; #(2*htp); // Sample(336)
        x =                0; #(2*htp); // Sample(337)
        x =              183; #(2*htp); // Sample(338)
        x =              290; #(2*htp); // Sample(339)
        x =              277; #(2*htp); // Sample(340)
        x =              150; #(2*htp); // Sample(341)
        x =              -39; #(2*htp); // Sample(342)
*/
        $finish;
    end
endmodule
