`timescale 1ns / 1ps

module testbench;

    // Inputs
    reg clk, reset;
    reg signed [31:0] x;
    wire signed [31:0] yw1;
    wire signed [31:0] y;
    // Instantiate the Unit Under Test (UUT)
    iir_order2 DUT(
      .clk(clk),
      .rst(reset),
      .x(x),
      .yw1(yw1),
      .y(y)
    );

    // Generate clock with 100ns period
    initial clk = 0;
    always #5 clk = ~clk;
    
    always @(posedge(clk)) begin
//      $display("time = %.0f,\t x = %.0f,\t w1->w2 = %.0f --> %.0f", $time, x, yw1, y);
      $display("%.0f,%.0f", x, y);
    end
    

    initial begin
        x = 32'd0;
        reset = 1;
        clk = 0;
        clk = 1;
        #10;
        reset = 0;
        #20;

        x =               25; #10; // Sample(1)
        x =               10; #10; // Sample(1)
        x =               25; #10; // Sample(1)
        x =               10; #10; // Sample(1)
        x =               67; #10; // Sample(1)
        x =              -56; #10; // Sample(2)
        x =               19; #10; // Sample(3)
        x =               28; #10; // Sample(4)
        x =              160; #10; // Sample(5)
        x =               39; #10; // Sample(6)
        x =              142; #10; // Sample(7)
        x =              151; #10; // Sample(8)
        x =              117; #10; // Sample(9)
        x =              294; #10; // Sample(10)
        x =              199; #10; // Sample(11)
        x =              363; #10; // Sample(12)
        x =              100; #10; // Sample(13)
        x =              525; #10; // Sample(14)
        x =               78; #10; // Sample(15)
        x =              195; #10; // Sample(16)
        x =              -19; #10; // Sample(17)
        x =              147; #10; // Sample(18)
        x =              515; #10; // Sample(19)
        x =              373; #10; // Sample(20)
        x =              110; #10; // Sample(21)
        x =              389; #10; // Sample(22)
        x =              161; #10; // Sample(23)
        x =              -98; #10; // Sample(24)
        x =              198; #10; // Sample(25)
        x =              673; #10; // Sample(26)
        x =              338; #10; // Sample(27)
        x =              -79; #10; // Sample(28)
        x =              424; #10; // Sample(29)
        x =              653; #10; // Sample(30)
        x =              269; #10; // Sample(31)
        x =              241; #10; // Sample(32)
        x =              374; #10; // Sample(33)
        x =               92; #10; // Sample(34)
        x =              296; #10; // Sample(35)
        x =              707; #10; // Sample(36)
        x =               46; #10; // Sample(37)
        x =              212; #10; // Sample(38)
        x =              262; #10; // Sample(39)
        x =              251; #10; // Sample(40)
        x =              315; #10; // Sample(41)
        x =               94; #10; // Sample(42)
        x =              -26; #10; // Sample(43)
        x =               84; #10; // Sample(44)
        x =             -286; #10; // Sample(45)
        x =               18; #10; // Sample(46)
        x =              459; #10; // Sample(47)
        x =              -86; #10; // Sample(48)
        x =               70; #10; // Sample(49)
        x =               77; #10; // Sample(50)
        x =               38; #10; // Sample(51)
        x =              -44; #10; // Sample(52)
        x =             -200; #10; // Sample(53)
        x =              -27; #10; // Sample(54)
        x =              -67; #10; // Sample(55)
        x =             -100; #10; // Sample(56)
        x =              -33; #10; // Sample(57)
        x =             -199; #10; // Sample(58)
        x =             -407; #10; // Sample(59)
        x =             -343; #10; // Sample(60)
        x =              -78; #10; // Sample(61)
        x =              -28; #10; // Sample(62)
        x =             -358; #10; // Sample(63)
        x =             -503; #10; // Sample(64)
        x =             -454; #10; // Sample(65)
        x =              -75; #10; // Sample(66)
        x =             -101; #10; // Sample(67)
        x =             -133; #10; // Sample(68)
        x =             -103; #10; // Sample(69)
        x =             -299; #10; // Sample(70)
        x =             -267; #10; // Sample(71)
        x =             -161; #10; // Sample(72)
        x =             -123; #10; // Sample(73)
        x =              191; #10; // Sample(74)
        x =             -482; #10; // Sample(75)
        x =             -272; #10; // Sample(76)
        x =             -206; #10; // Sample(77)
        x =             -506; #10; // Sample(78)
        x =             -562; #10; // Sample(79)
        x =             -238; #10; // Sample(80)
        x =             -396; #10; // Sample(81)
        x =             -249; #10; // Sample(82)
        x =             -421; #10; // Sample(83)
        x =             -245; #10; // Sample(84)
        x =             -193; #10; // Sample(85)
        x =             -624; #10; // Sample(86)
        x =              -37; #10; // Sample(87)
        x =             -554; #10; // Sample(88)
        x =             -101; #10; // Sample(89)
        x =             -129; #10; // Sample(90)
        x =              -70; #10; // Sample(91)
        x =              197; #10; // Sample(92)
        x =             -374; #10; // Sample(93)
        x =             -191; #10; // Sample(94)
        x =             -186; #10; // Sample(95)
        x =              278; #10; // Sample(96)
        x =              253; #10; // Sample(97)
        x =              156; #10; // Sample(98)
        x =             -260; #10; // Sample(99)
        x =              -30; #10; // Sample(100)
        x =              179; #10; // Sample(101)
        x =              164; #10; // Sample(102)
        x =              -10; #10; // Sample(103)
        x =              423; #10; // Sample(104)
        x =               39; #10; // Sample(105)
        x =              241; #10; // Sample(106)
        x =              568; #10; // Sample(107)
        x =              532; #10; // Sample(108)
        x =              174; #10; // Sample(109)
        x =              371; #10; // Sample(110)
        x =              562; #10; // Sample(111)
        x =               66; #10; // Sample(112)
        x =              445; #10; // Sample(113)
        x =              628; #10; // Sample(114)
        x =              471; #10; // Sample(115)
        x =              522; #10; // Sample(116)
        x =              290; #10; // Sample(117)
        x =               47; #10; // Sample(118)
        x =              157; #10; // Sample(119)
        x =              597; #10; // Sample(120)
        x =              314; #10; // Sample(121)
        x =              458; #10; // Sample(122)
        x =              102; #10; // Sample(123)
        x =              -47; #10; // Sample(124)
        x =             -105; #10; // Sample(125)
        x =              338; #10; // Sample(126)
        x =             -133; #10; // Sample(127)
        x =              543; #10; // Sample(128)
        x =              479; #10; // Sample(129)
        x =              307; #10; // Sample(130)
        x =              435; #10; // Sample(131)
        x =              206; #10; // Sample(132)
        x =             -133; #10; // Sample(133)
        x =              174; #10; // Sample(134)
        x =               55; #10; // Sample(135)
        x =              405; #10; // Sample(136)
        x =              216; #10; // Sample(137)
        x =              211; #10; // Sample(138)
        x =               45; #10; // Sample(139)
        x =              -72; #10; // Sample(140)
        x =              131; #10; // Sample(141)
        x =              -23; #10; // Sample(142)
        x =              301; #10; // Sample(143)
        x =              -49; #10; // Sample(144)
        x =             -150; #10; // Sample(145)
        x =              -61; #10; // Sample(146)
        x =              165; #10; // Sample(147)
        x =             -166; #10; // Sample(148)
        x =              -96; #10; // Sample(149)
        x =             -374; #10; // Sample(150)
        x =              -92; #10; // Sample(151)
        x =             -205; #10; // Sample(152)
        x =             -234; #10; // Sample(153)
        x =             -140; #10; // Sample(154)
        x =             -178; #10; // Sample(155)
        x =             -198; #10; // Sample(156)
        x =              354; #10; // Sample(157)
        x =              -29; #10; // Sample(158)
        x =               80; #10; // Sample(159)
        x =               65; #10; // Sample(160)
        x =             -314; #10; // Sample(161)
        x =             -361; #10; // Sample(162)
        x =             -591; #10; // Sample(163)
        x =             -467; #10; // Sample(164)
        x =             -344; #10; // Sample(165)
        x =             -311; #10; // Sample(166)
        x =             -236; #10; // Sample(167)
        x =             -270; #10; // Sample(168)
        x =             -525; #10; // Sample(169)
        x =             -361; #10; // Sample(170)
        x =               30; #10; // Sample(171)
        x =             -351; #10; // Sample(172)
        x =             -464; #10; // Sample(173)
        x =             -332; #10; // Sample(174)
        x =             -214; #10; // Sample(175)
        x =             -342; #10; // Sample(176)
        x =             -341; #10; // Sample(177)
        x =             -314; #10; // Sample(178)
        x =              -13; #10; // Sample(179)
        x =              -67; #10; // Sample(180)
        x =             -354; #10; // Sample(181)
        x =             -339; #10; // Sample(182)
        x =             -512; #10; // Sample(183)
        x =               46; #10; // Sample(184)
        x =             -170; #10; // Sample(185)
        x =             -179; #10; // Sample(186)
        x =              -81; #10; // Sample(187)
        x =             -342; #10; // Sample(188)
        x =             -252; #10; // Sample(189)
        x =              -24; #10; // Sample(190)
        x =             -100; #10; // Sample(191)
        x =             -409; #10; // Sample(192)
        x =             -146; #10; // Sample(193)
        x =               70; #10; // Sample(194)
        x =              242; #10; // Sample(195)
        x =               76; #10; // Sample(196)
        x =              105; #10; // Sample(197)
        x =                5; #10; // Sample(198)
        x =              155; #10; // Sample(199)
        x =              236; #10; // Sample(200)
        x =              -21; #10; // Sample(201)
        x =              366; #10; // Sample(202)
        x =             -132; #10; // Sample(203)
        x =              189; #10; // Sample(204)
        x =              168; #10; // Sample(205)
        x =              538; #10; // Sample(206)
        x =              179; #10; // Sample(207)
        x =              861; #10; // Sample(208)
        x =              208; #10; // Sample(209)
        x =              133; #10; // Sample(210)
        x =              718; #10; // Sample(211)
        x =              280; #10; // Sample(212)
        x =              241; #10; // Sample(213)
        x =              322; #10; // Sample(214)
        x =              107; #10; // Sample(215)
        x =               22; #10; // Sample(216)
        x =              178; #10; // Sample(217)
        x =              312; #10; // Sample(218)
        x =              514; #10; // Sample(219)
        x =              524; #10; // Sample(220)
        x =              381; #10; // Sample(221)
        x =              511; #10; // Sample(222)
        x =              775; #10; // Sample(223)
        x =              393; #10; // Sample(224)
        x =              443; #10; // Sample(225)
        x =              192; #10; // Sample(226)
        x =              466; #10; // Sample(227)
        x =               12; #10; // Sample(228)
        x =              149; #10; // Sample(229)
        x =               35; #10; // Sample(230)
        x =               77; #10; // Sample(231)
        x =              545; #10; // Sample(232)
        x =              111; #10; // Sample(233)
        x =               52; #10; // Sample(234)
        x =              311; #10; // Sample(235)
        x =               36; #10; // Sample(236)
        x =              139; #10; // Sample(237)
        x =              164; #10; // Sample(238)
        x =             -126; #10; // Sample(239)
        x =              -47; #10; // Sample(240)
        x =              365; #10; // Sample(241)
        x =                6; #10; // Sample(242)
        x =              133; #10; // Sample(243)
        x =              184; #10; // Sample(244)
        x =               32; #10; // Sample(245)
        x =              -72; #10; // Sample(246)
        x =              129; #10; // Sample(247)
        x =             -372; #10; // Sample(248)
        x =               80; #10; // Sample(249)
        x =             -567; #10; // Sample(250)
        x =             -423; #10; // Sample(251)
        x =             -279; #10; // Sample(252)
        x =             -228; #10; // Sample(253)
        x =             -536; #10; // Sample(254)
        x =              -90; #10; // Sample(255)
        x =             -264; #10; // Sample(256)
        x =             -469; #10; // Sample(257)
        x =             -496; #10; // Sample(258)
        x =             -460; #10; // Sample(259)
        x =             -443; #10; // Sample(260)
        x =             -314; #10; // Sample(261)
        x =             -304; #10; // Sample(262)
        x =             -408; #10; // Sample(263)
        x =             -315; #10; // Sample(264)
        x =             -423; #10; // Sample(265)
        x =             -265; #10; // Sample(266)
        x =               -2; #10; // Sample(267)
        x =             -130; #10; // Sample(268)
        x =             -368; #10; // Sample(269)
        x =             -256; #10; // Sample(270)
        x =             -307; #10; // Sample(271)
        x =             -350; #10; // Sample(272)
        x =             -320; #10; // Sample(273)
        x =              -38; #10; // Sample(274)
        x =             -342; #10; // Sample(275)
        x =             -190; #10; // Sample(276)
        x =              -95; #10; // Sample(277)
        x =             -395; #10; // Sample(278)
        x =             -470; #10; // Sample(279)
        x =              -21; #10; // Sample(280)
        x =              -77; #10; // Sample(281)
        x =             -235; #10; // Sample(282)
        x =              100; #10; // Sample(283)
        x =              -36; #10; // Sample(284)
        x =             -155; #10; // Sample(285)
        x =             -143; #10; // Sample(286)
        x =             -134; #10; // Sample(287)
        x =             -228; #10; // Sample(288)
        x =              519; #10; // Sample(289)
        x =             -412; #10; // Sample(290)
        x =               91; #10; // Sample(291)
        x =               60; #10; // Sample(292)
        x =             -166; #10; // Sample(293)
        x =               68; #10; // Sample(294)
        x =              189; #10; // Sample(295)
        x =              328; #10; // Sample(296)
        x =              171; #10; // Sample(297)
        x =              278; #10; // Sample(298)
        x =              516; #10; // Sample(299)
        x =              177; #10; // Sample(300)
        x =              103; #10; // Sample(301)
        x =              -46; #10; // Sample(302)
        x =              399; #10; // Sample(303)
        x =              152; #10; // Sample(304)
        x =              530; #10; // Sample(305)
        x =              283; #10; // Sample(306)
        x =              251; #10; // Sample(307)
        x =              177; #10; // Sample(308)
        x =              192; #10; // Sample(309)
        x =               54; #10; // Sample(310)
        x =              411; #10; // Sample(311)
        x =              219; #10; // Sample(312)
        x =              421; #10; // Sample(313)
        x =              -22; #10; // Sample(314)
        x =              362; #10; // Sample(315)
        x =              120; #10; // Sample(316)
        x =               -7; #10; // Sample(317)
        x =              239; #10; // Sample(318)
        x =              394; #10; // Sample(319)
        x =              465; #10; // Sample(320)
        x =              494; #10; // Sample(321)
        x =              177; #10; // Sample(322)
        x =               56; #10; // Sample(323)
        x =              802; #10; // Sample(324)
        x =              108; #10; // Sample(325)
        x =               64; #10; // Sample(326)
        x =              273; #10; // Sample(327)
        x =              -37; #10; // Sample(328)
        x =               24; #10; // Sample(329)
        x =             -156; #10; // Sample(330)
        x =               77; #10; // Sample(331)
        x =             -117; #10; // Sample(332)
        x =              152; #10; // Sample(333)
        x =               95; #10; // Sample(334)
        x =              -97; #10; // Sample(335)
        x =              -53; #10; // Sample(336)
        x =             -108; #10; // Sample(337)
        x =               12; #10; // Sample(338)
        x =             -163; #10; // Sample(339)
        x =               -8; #10; // Sample(340)
        x =             -239; #10; // Sample(341)
        x =               15; #10; // Sample(342)
        x =             -146; #10; // Sample(343)
        x =             -521; #10; // Sample(344)
        x =             -114; #10; // Sample(345)
        x =               12; #10; // Sample(346)
        x =               56; #10; // Sample(347)
        x =             -155; #10; // Sample(348)
        x =               68; #10; // Sample(349)
        x =              -95; #10; // Sample(350)
        x =              160; #10; // Sample(351)
        x =             -199; #10; // Sample(352)
        x =             -169; #10; // Sample(353)
        x =             -187; #10; // Sample(354)
        x =             -172; #10; // Sample(355)
        x =             -127; #10; // Sample(356)
        x =              -89; #10; // Sample(357)
        x =             -480; #10; // Sample(358)
        x =             -542; #10; // Sample(359)
        x =              -47; #10; // Sample(360)
        x =             -117; #10; // Sample(361)
        x =             -459; #10; // Sample(362)
        x =             -306; #10; // Sample(363)
        x =               55; #10; // Sample(364)
        x =             -508; #10; // Sample(365)
        x =             -222; #10; // Sample(366)
        x =             -539; #10; // Sample(367)
        x =             -236; #10; // Sample(368)
        x =             -202; #10; // Sample(369)
        x =             -283; #10; // Sample(370)
        x =              -60; #10; // Sample(371)
        x =             -252; #10; // Sample(372)
        x =               12; #10; // Sample(373)
        x =                9; #10; // Sample(374)
        x =             -235; #10; // Sample(375)
        x =             -118; #10; // Sample(376)
        x =             -110; #10; // Sample(377)
        x =               50; #10; // Sample(378)
        x =              120; #10; // Sample(379)
        x =               54; #10; // Sample(380)
        x =              -73; #10; // Sample(381)
        x =             -227; #10; // Sample(382)
        x =             -282; #10; // Sample(383)
        x =              188; #10; // Sample(384)
        x =              377; #10; // Sample(385)
        x =               71; #10; // Sample(386)
        x =               26; #10; // Sample(387)
        x =              236; #10; // Sample(388)
        x =             -239; #10; // Sample(389)
        x =               47; #10; // Sample(390)
        x =             -262; #10; // Sample(391)
        x =              214; #10; // Sample(392)
        x =              156; #10; // Sample(393)
        x =              229; #10; // Sample(394)
        x =              102; #10; // Sample(395)
        x =             -154; #10; // Sample(396)
        x =              400; #10; // Sample(397)
        x =              103; #10; // Sample(398)
        x =              272; #10; // Sample(399)
        x =              429; #10; // Sample(400)
        x =              368; #10; // Sample(401)
        x =              113; #10; // Sample(402)
        x =              228; #10; // Sample(403)
        x =              243; #10; // Sample(404)
        x =              477; #10; // Sample(405)
        x =              537; #10; // Sample(406)
        x =               97; #10; // Sample(407)
        x =              107; #10; // Sample(408)
        x =              325; #10; // Sample(409)
        x =              299; #10; // Sample(410)
        x =              335; #10; // Sample(411)
        x =               96; #10; // Sample(412)
        x =               37; #10; // Sample(413)
        x =              269; #10; // Sample(414)
        x =              511; #10; // Sample(415)
        x =              389; #10; // Sample(416)
        x =              238; #10; // Sample(417)
        x =              177; #10; // Sample(418)
        x =               26; #10; // Sample(419)
        x =              396; #10; // Sample(420)
        x =              374; #10; // Sample(421)
        x =              167; #10; // Sample(422)
        x =              256; #10; // Sample(423)
        x =              219; #10; // Sample(424)
        x =              325; #10; // Sample(425)
        x =              443; #10; // Sample(426)
        x =             -217; #10; // Sample(427)
        x =               38; #10; // Sample(428)
        x =               63; #10; // Sample(429)
        x =             -182; #10; // Sample(430)
        x =              -16; #10; // Sample(431)
        x =              174; #10; // Sample(432)
        x =             -143; #10; // Sample(433)
        x =             -417; #10; // Sample(434)
        x =             -232; #10; // Sample(435)
        x =               -5; #10; // Sample(436)
        x =             -222; #10; // Sample(437)
        x =               83; #10; // Sample(438)
        x =             -220; #10; // Sample(439)
        x =              -89; #10; // Sample(440)
        x =             -263; #10; // Sample(441)
        x =              -48; #10; // Sample(442)
        x =             -493; #10; // Sample(443)
        x =              112; #10; // Sample(444)
        x =             -253; #10; // Sample(445)
        x =             -252; #10; // Sample(446)
        x =             -507; #10; // Sample(447)
        x =             -249; #10; // Sample(448)
        x =             -273; #10; // Sample(449)
        x =             -497; #10; // Sample(450)
        x =             -164; #10; // Sample(451)
        x =               96; #10; // Sample(452)
        x =              -65; #10; // Sample(453)
        x =             -306; #10; // Sample(454)
        x =             -192; #10; // Sample(455)
        x =             -259; #10; // Sample(456)
        x =             -221; #10; // Sample(457)
        x =             -689; #10; // Sample(458)
        x =             -468; #10; // Sample(459)
        x =             -348; #10; // Sample(460)
        x =             -170; #10; // Sample(461)
        x =             -215; #10; // Sample(462)
        x =             -296; #10; // Sample(463)
        x =             -677; #10; // Sample(464)
        x =             -529; #10; // Sample(465)
        x =                4; #10; // Sample(466)
        x =             -212; #10; // Sample(467)
        x =             -223; #10; // Sample(468)
        x =             -276; #10; // Sample(469)
        x =              351; #10; // Sample(470)
        x =             -312; #10; // Sample(471)
        x =             -194; #10; // Sample(472)
        x =              -49; #10; // Sample(473)
        x =              117; #10; // Sample(474)
        x =             -140; #10; // Sample(475)
        x =               87; #10; // Sample(476)
        x =              110; #10; // Sample(477)
        x =              -10; #10; // Sample(478)
        x =             -287; #10; // Sample(479)
        x =              132; #10; // Sample(480)
        x =               20; #10; // Sample(481)
        x =              313; #10; // Sample(482)
        x =             -119; #10; // Sample(483)
        x =               58; #10; // Sample(484)
        x =              -17; #10; // Sample(485)
        x =             -251; #10; // Sample(486)
        x =              -83; #10; // Sample(487)
        x =             -236; #10; // Sample(488)
        x =              469; #10; // Sample(489)
        x =              213; #10; // Sample(490)
        x =              296; #10; // Sample(491)
        x =              237; #10; // Sample(492)
        x =              423; #10; // Sample(493)
        x =              512; #10; // Sample(494)
        x =              162; #10; // Sample(495)
        x =               67; #10; // Sample(496)
        x =              469; #10; // Sample(497)
        x =              693; #10; // Sample(498)
        x =              236; #10; // Sample(499)
        x =              141; #10; // Sample(500)
        x =                0; #10; // Sample(1)
        x =              183; #10; // Sample(2)
        x =              290; #10; // Sample(3)
        x =              277; #10; // Sample(4)
        x =              150; #10; // Sample(5)
        x =              -39; #10; // Sample(6)
        x =             -212; #10; // Sample(7)
        x =             -297; #10; // Sample(8)
        x =             -260; #10; // Sample(9)
        x =             -115; #10; // Sample(10)
        x =               78; #10; // Sample(11)
        x =              238; #10; // Sample(12)
        x =              300; #10; // Sample(13)
        x =              238; #10; // Sample(14)
        x =               78; #10; // Sample(15)
        x =             -115; #10; // Sample(16)
        x =             -260; #10; // Sample(17)
        x =             -297; #10; // Sample(18)
        x =             -212; #10; // Sample(19)
        x =              -39; #10; // Sample(20)
        x =              150; #10; // Sample(21)
        x =              277; #10; // Sample(22)
        x =              290; #10; // Sample(23)
        x =              183; #10; // Sample(24)
        x =                0; #10; // Sample(25)
        x =             -183; #10; // Sample(26)
        x =             -290; #10; // Sample(27)
        x =             -277; #10; // Sample(28)
        x =             -150; #10; // Sample(29)
        x =               39; #10; // Sample(30)
        x =              212; #10; // Sample(31)
        x =              297; #10; // Sample(32)
        x =              260; #10; // Sample(33)
        x =              115; #10; // Sample(34)
        x =              -78; #10; // Sample(35)
        x =             -238; #10; // Sample(36)
        x =             -300; #10; // Sample(37)
        x =             -238; #10; // Sample(38)
        x =              -78; #10; // Sample(39)
        x =              115; #10; // Sample(40)
        x =              260; #10; // Sample(41)
        x =              297; #10; // Sample(42)
        x =              212; #10; // Sample(43)
        x =               39; #10; // Sample(44)
        x =             -150; #10; // Sample(45)
        x =             -277; #10; // Sample(46)
        x =             -290; #10; // Sample(47)
        x =             -183; #10; // Sample(48)
        x =               -0; #10; // Sample(49)
        x =              183; #10; // Sample(50)
        x =              290; #10; // Sample(51)
        x =              277; #10; // Sample(52)

/*
        x =              150; #10; // Sample(53)
        x =              -39; #10; // Sample(54)
        x =             -212; #10; // Sample(55)
        x =             -297; #10; // Sample(56)
        x =             -260; #10; // Sample(57)
        x =             -115; #10; // Sample(58)
        x =               78; #10; // Sample(59)
        x =              238; #10; // Sample(60)
        x =              300; #10; // Sample(61)
        x =              238; #10; // Sample(62)
        x =               78; #10; // Sample(63)
        x =             -115; #10; // Sample(64)
        x =             -260; #10; // Sample(65)
        x =             -297; #10; // Sample(66)
        x =             -212; #10; // Sample(67)
        x =              -39; #10; // Sample(68)
        x =              150; #10; // Sample(69)
        x =              277; #10; // Sample(70)
        x =              290; #10; // Sample(71)
        x =              183; #10; // Sample(72)
        x =               -0; #10; // Sample(73)
        x =             -183; #10; // Sample(74)
        x =             -290; #10; // Sample(75)
        x =             -277; #10; // Sample(76)
        x =             -150; #10; // Sample(77)
        x =               39; #10; // Sample(78)
        x =              212; #10; // Sample(79)
        x =              297; #10; // Sample(80)
        x =              260; #10; // Sample(81)
        x =              115; #10; // Sample(82)
        x =              -78; #10; // Sample(83)
        x =             -238; #10; // Sample(84)
        x =             -300; #10; // Sample(85)
        x =             -238; #10; // Sample(86)
        x =              -78; #10; // Sample(87)
        x =              115; #10; // Sample(88)
        x =              260; #10; // Sample(89)
        x =              297; #10; // Sample(90)
        x =              212; #10; // Sample(91)
        x =               39; #10; // Sample(92)
        x =             -150; #10; // Sample(93)
        x =             -277; #10; // Sample(94)
        x =             -290; #10; // Sample(95)
        x =             -183; #10; // Sample(96)
        x =               -0; #10; // Sample(97)
        x =              183; #10; // Sample(98)
        x =              290; #10; // Sample(99)
        x =              277; #10; // Sample(100)
        x =              150; #10; // Sample(101)
        x =              -39; #10; // Sample(102)
        x =             -212; #10; // Sample(103)
        x =             -297; #10; // Sample(104)
        x =             -260; #10; // Sample(105)
        x =             -115; #10; // Sample(106)
        x =               78; #10; // Sample(107)
        x =              238; #10; // Sample(108)
        x =              300; #10; // Sample(109)
        x =              238; #10; // Sample(110)
        x =               78; #10; // Sample(111)
        x =             -115; #10; // Sample(112)
        x =             -260; #10; // Sample(113)
        x =             -297; #10; // Sample(114)
        x =             -212; #10; // Sample(115)
        x =              -39; #10; // Sample(116)
        x =              150; #10; // Sample(117)
        x =              277; #10; // Sample(118)
        x =              290; #10; // Sample(119)
        x =              183; #10; // Sample(120)
        x =               -0; #10; // Sample(121)
        x =             -183; #10; // Sample(122)
        x =             -290; #10; // Sample(123)
        x =             -277; #10; // Sample(124)
        x =             -150; #10; // Sample(125)
        x =               39; #10; // Sample(126)
        x =              212; #10; // Sample(127)
        x =              297; #10; // Sample(128)
        x =              260; #10; // Sample(129)
        x =              115; #10; // Sample(130)
        x =              -78; #10; // Sample(131)
        x =             -238; #10; // Sample(132)
        x =             -300; #10; // Sample(133)
        x =             -238; #10; // Sample(134)
        x =              -78; #10; // Sample(135)
        x =              115; #10; // Sample(136)
        x =              260; #10; // Sample(137)
        x =              297; #10; // Sample(138)
        x =              212; #10; // Sample(139)
        x =               39; #10; // Sample(140)
        x =             -150; #10; // Sample(141)
        x =             -277; #10; // Sample(142)
        x =             -290; #10; // Sample(143)
        x =             -183; #10; // Sample(144)
        x =                0; #10; // Sample(145)
        x =              183; #10; // Sample(146)
        x =              290; #10; // Sample(147)
        x =              277; #10; // Sample(148)
        x =              150; #10; // Sample(149)
        x =              -39; #10; // Sample(150)
        x =             -212; #10; // Sample(151)
        x =             -297; #10; // Sample(152)
        x =             -260; #10; // Sample(153)
        x =             -115; #10; // Sample(154)
        x =               78; #10; // Sample(155)
        x =              238; #10; // Sample(156)
        x =              300; #10; // Sample(157)
        x =              238; #10; // Sample(158)
        x =               78; #10; // Sample(159)
        x =             -115; #10; // Sample(160)
        x =             -260; #10; // Sample(161)
        x =             -297; #10; // Sample(162)
        x =             -212; #10; // Sample(163)
        x =              -39; #10; // Sample(164)
        x =              150; #10; // Sample(165)
        x =              277; #10; // Sample(166)
        x =              290; #10; // Sample(167)
        x =              183; #10; // Sample(168)
        x =               -0; #10; // Sample(169)
        x =             -183; #10; // Sample(170)
        x =             -290; #10; // Sample(171)
        x =             -277; #10; // Sample(172)
        x =             -150; #10; // Sample(173)
        x =               39; #10; // Sample(174)
        x =              212; #10; // Sample(175)
        x =              297; #10; // Sample(176)
        x =              260; #10; // Sample(177)
        x =              115; #10; // Sample(178)
        x =              -78; #10; // Sample(179)
        x =             -238; #10; // Sample(180)
        x =             -300; #10; // Sample(181)
        x =             -238; #10; // Sample(182)
        x =              -78; #10; // Sample(183)
        x =              115; #10; // Sample(184)
        x =              260; #10; // Sample(185)
        x =              297; #10; // Sample(186)
        x =              212; #10; // Sample(187)
        x =               39; #10; // Sample(188)
        x =             -150; #10; // Sample(189)
        x =             -277; #10; // Sample(190)
        x =             -290; #10; // Sample(191)
        x =             -183; #10; // Sample(192)
        x =               -0; #10; // Sample(193)
        x =              183; #10; // Sample(194)
        x =              290; #10; // Sample(195)
        x =              277; #10; // Sample(196)
        x =              150; #10; // Sample(197)
        x =              -39; #10; // Sample(198)
        x =             -212; #10; // Sample(199)
        x =             -297; #10; // Sample(200)
        x =             -260; #10; // Sample(201)
        x =             -115; #10; // Sample(202)
        x =               78; #10; // Sample(203)
        x =              238; #10; // Sample(204)
        x =              300; #10; // Sample(205)
        x =              238; #10; // Sample(206)
        x =               78; #10; // Sample(207)
        x =             -115; #10; // Sample(208)
        x =             -260; #10; // Sample(209)
        x =             -297; #10; // Sample(210)
        x =             -212; #10; // Sample(211)
        x =              -39; #10; // Sample(212)
        x =              150; #10; // Sample(213)
        x =              277; #10; // Sample(214)
        x =              290; #10; // Sample(215)
        x =              183; #10; // Sample(216)
        x =                0; #10; // Sample(217)
        x =             -183; #10; // Sample(218)
        x =             -290; #10; // Sample(219)
        x =             -277; #10; // Sample(220)
        x =             -150; #10; // Sample(221)
        x =               39; #10; // Sample(222)
        x =              212; #10; // Sample(223)
        x =              297; #10; // Sample(224)
        x =              260; #10; // Sample(225)
        x =              115; #10; // Sample(226)
        x =              -78; #10; // Sample(227)
        x =             -238; #10; // Sample(228)
        x =             -300; #10; // Sample(229)
        x =             -238; #10; // Sample(230)
        x =              -78; #10; // Sample(231)
        x =              115; #10; // Sample(232)
        x =              260; #10; // Sample(233)
        x =              297; #10; // Sample(234)
        x =              212; #10; // Sample(235)
        x =               39; #10; // Sample(236)
        x =             -150; #10; // Sample(237)
        x =             -277; #10; // Sample(238)
        x =             -290; #10; // Sample(239)
        x =             -183; #10; // Sample(240)
        x =                0; #10; // Sample(241)
        x =              183; #10; // Sample(242)
        x =              290; #10; // Sample(243)
        x =              277; #10; // Sample(244)
        x =              150; #10; // Sample(245)
        x =              -39; #10; // Sample(246)
        x =             -212; #10; // Sample(247)
        x =             -297; #10; // Sample(248)
        x =             -260; #10; // Sample(249)
        x =             -115; #10; // Sample(250)
        x =               78; #10; // Sample(251)
        x =              238; #10; // Sample(252)
        x =              300; #10; // Sample(253)
        x =              238; #10; // Sample(254)
        x =               78; #10; // Sample(255)
        x =             -115; #10; // Sample(256)
        x =             -260; #10; // Sample(257)
        x =             -297; #10; // Sample(258)
        x =             -212; #10; // Sample(259)
        x =              -39; #10; // Sample(260)
        x =              150; #10; // Sample(261)
        x =              277; #10; // Sample(262)
        x =              290; #10; // Sample(263)
        x =              183; #10; // Sample(264)
        x =               -0; #10; // Sample(265)
        x =             -183; #10; // Sample(266)
        x =             -290; #10; // Sample(267)
        x =             -277; #10; // Sample(268)
        x =             -150; #10; // Sample(269)
        x =               39; #10; // Sample(270)
        x =              212; #10; // Sample(271)
        x =              297; #10; // Sample(272)
        x =              260; #10; // Sample(273)
        x =              115; #10; // Sample(274)
        x =              -78; #10; // Sample(275)
        x =             -238; #10; // Sample(276)
        x =             -300; #10; // Sample(277)
        x =             -238; #10; // Sample(278)
        x =              -78; #10; // Sample(279)
        x =              115; #10; // Sample(280)
        x =              260; #10; // Sample(281)
        x =              297; #10; // Sample(282)
        x =              212; #10; // Sample(283)
        x =               39; #10; // Sample(284)
        x =             -150; #10; // Sample(285)
        x =             -277; #10; // Sample(286)
        x =             -290; #10; // Sample(287)
        x =             -183; #10; // Sample(288)
        x =                0; #10; // Sample(289)
        x =              183; #10; // Sample(290)
        x =              290; #10; // Sample(291)
        x =              277; #10; // Sample(292)
        x =              150; #10; // Sample(293)
        x =              -39; #10; // Sample(294)
        x =             -212; #10; // Sample(295)
        x =             -297; #10; // Sample(296)
        x =             -260; #10; // Sample(297)
        x =             -115; #10; // Sample(298)
        x =               78; #10; // Sample(299)
        x =              238; #10; // Sample(300)
        x =              300; #10; // Sample(301)
        x =              238; #10; // Sample(302)
        x =               78; #10; // Sample(303)
        x =             -115; #10; // Sample(304)
        x =             -260; #10; // Sample(305)
        x =             -297; #10; // Sample(306)
        x =             -212; #10; // Sample(307)
        x =              -39; #10; // Sample(308)
        x =              150; #10; // Sample(309)
        x =              277; #10; // Sample(310)
        x =              290; #10; // Sample(311)
        x =              183; #10; // Sample(312)
        x =               -0; #10; // Sample(313)
        x =             -183; #10; // Sample(314)
        x =             -290; #10; // Sample(315)
        x =             -277; #10; // Sample(316)
        x =             -150; #10; // Sample(317)
        x =               39; #10; // Sample(318)
        x =              212; #10; // Sample(319)
        x =              297; #10; // Sample(320)
        x =              260; #10; // Sample(321)
        x =              115; #10; // Sample(322)
        x =              -78; #10; // Sample(323)
        x =             -238; #10; // Sample(324)
        x =             -300; #10; // Sample(325)
        x =             -238; #10; // Sample(326)
        x =              -78; #10; // Sample(327)
        x =              115; #10; // Sample(328)
        x =              260; #10; // Sample(329)
        x =              297; #10; // Sample(330)
        x =              212; #10; // Sample(331)
        x =               39; #10; // Sample(332)
        x =             -150; #10; // Sample(333)
        x =             -277; #10; // Sample(334)
        x =             -290; #10; // Sample(335)
        x =             -183; #10; // Sample(336)
        x =                0; #10; // Sample(337)
        x =              183; #10; // Sample(338)
        x =              290; #10; // Sample(339)
        x =              277; #10; // Sample(340)
        x =              150; #10; // Sample(341)
        x =              -39; #10; // Sample(342)
*/
        $finish;
    end
endmodule
