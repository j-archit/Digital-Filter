`timescale 1ns / 1ps

module testbench;

    // Inputs
    reg clk, reset;
    reg signed [31:0] x;
    wire signed [31:0] t;
    wire signed [31:0] t2;
    wire signed [31:0] t3;
    wire signed [31:0] y;

    // Instantiate the Unit Under Test (UUT)
    iir_order2 DUT1(
      .clk(clk),
      .rst(reset),
      .x(x),
      .y(t)
    );
    iir_order2 DUT2(
      .clk(clk),
      .rst(reset),
      .x(t),
      .y(y)
    );

    // Generate clock with 100ns period
    initial clk = 0;
    always #25 clk = ~clk;
    
    always @(posedge(clk)) begin
//      $display("time = %.0f,\t x = %.0f,\t w2 = %.0f", $time, x, y);
      $display("%.0f,%.0f", x, y);
    end
    

    initial begin
        x = 32'd0;
        reset = 1;
        clk = 0;
        clk = 1;
        #10;
        reset = 0;
        #20;

        x =               25; #50; // Sample(1)
        x =               10; #50; // Sample(1)
        x =               25; #50; // Sample(1)
        x =               10; #50; // Sample(1)
        x =               67; #50; // Sample(1)
        x =              -56; #50; // Sample(2)
        x =               19; #50; // Sample(3)
        x =               28; #50; // Sample(4)
        x =              160; #50; // Sample(5)
        x =               39; #50; // Sample(6)
        x =              142; #50; // Sample(7)
        x =              151; #50; // Sample(8)
        x =              117; #50; // Sample(9)
        x =              294; #50; // Sample(10)
        x =              199; #50; // Sample(11)
        x =              363; #50; // Sample(12)
        x =              100; #50; // Sample(13)
        x =              525; #50; // Sample(14)
        x =               78; #50; // Sample(15)
        x =              195; #50; // Sample(16)
        x =              -19; #50; // Sample(17)
        x =              147; #50; // Sample(18)
        x =              515; #50; // Sample(19)
        x =              373; #50; // Sample(20)
        x =              110; #50; // Sample(21)
        x =              389; #50; // Sample(22)
        x =              161; #50; // Sample(23)
        x =              -98; #50; // Sample(24)
        x =              198; #50; // Sample(25)
        x =              673; #50; // Sample(26)
        x =              338; #50; // Sample(27)
        x =              -79; #50; // Sample(28)
        x =              424; #50; // Sample(29)
        x =              653; #50; // Sample(30)
        x =              269; #50; // Sample(31)
        x =              241; #50; // Sample(32)
        x =              374; #50; // Sample(33)
        x =               92; #50; // Sample(34)
        x =              296; #50; // Sample(35)
        x =              707; #50; // Sample(36)
        x =               46; #50; // Sample(37)
        x =              212; #50; // Sample(38)
        x =              262; #50; // Sample(39)
        x =              251; #50; // Sample(40)
        x =              315; #50; // Sample(41)
        x =               94; #50; // Sample(42)
        x =              -26; #50; // Sample(43)
        x =               84; #50; // Sample(44)
        x =             -286; #50; // Sample(45)
        x =               18; #50; // Sample(46)
        x =              459; #50; // Sample(47)
        x =              -86; #50; // Sample(48)
        x =               70; #50; // Sample(49)
        x =               77; #50; // Sample(50)
        x =               38; #50; // Sample(51)
        x =              -44; #50; // Sample(52)
        x =             -200; #50; // Sample(53)
        x =              -27; #50; // Sample(54)
        x =              -67; #50; // Sample(55)
        x =             -100; #50; // Sample(56)
        x =              -33; #50; // Sample(57)
        x =             -199; #50; // Sample(58)
        x =             -407; #50; // Sample(59)
        x =             -343; #50; // Sample(60)
        x =              -78; #50; // Sample(61)
        x =              -28; #50; // Sample(62)
        x =             -358; #50; // Sample(63)
        x =             -503; #50; // Sample(64)
        x =             -454; #50; // Sample(65)
        x =              -75; #50; // Sample(66)
        x =             -101; #50; // Sample(67)
        x =             -133; #50; // Sample(68)
        x =             -103; #50; // Sample(69)
        x =             -299; #50; // Sample(70)
        x =             -267; #50; // Sample(71)
        x =             -161; #50; // Sample(72)
        x =             -123; #50; // Sample(73)
        x =              191; #50; // Sample(74)
        x =             -482; #50; // Sample(75)
        x =             -272; #50; // Sample(76)
        x =             -206; #50; // Sample(77)
        x =             -506; #50; // Sample(78)
        x =             -562; #50; // Sample(79)
        x =             -238; #50; // Sample(80)
        x =             -396; #50; // Sample(81)
        x =             -249; #50; // Sample(82)
        x =             -421; #50; // Sample(83)
        x =             -245; #50; // Sample(84)
        x =             -193; #50; // Sample(85)
        x =             -624; #50; // Sample(86)
        x =              -37; #50; // Sample(87)
        x =             -554; #50; // Sample(88)
        x =             -101; #50; // Sample(89)
        x =             -129; #50; // Sample(90)
        x =              -70; #50; // Sample(91)
        x =              197; #50; // Sample(92)
        x =             -374; #50; // Sample(93)
        x =             -191; #50; // Sample(94)
        x =             -186; #50; // Sample(95)
        x =              278; #50; // Sample(96)
        x =              253; #50; // Sample(97)
        x =              156; #50; // Sample(98)
        x =             -260; #50; // Sample(99)
        x =              -30; #50; // Sample(100)
        x =              179; #50; // Sample(101)
        x =              164; #50; // Sample(102)
        x =              -10; #50; // Sample(103)
        x =              423; #50; // Sample(104)
        x =               39; #50; // Sample(105)
        x =              241; #50; // Sample(106)
        x =              568; #50; // Sample(107)
        x =              532; #50; // Sample(108)
        x =              174; #50; // Sample(109)
        x =              371; #50; // Sample(110)
        x =              562; #50; // Sample(111)
        x =               66; #50; // Sample(112)
        x =              445; #50; // Sample(113)
        x =              628; #50; // Sample(114)
        x =              471; #50; // Sample(115)
        x =              522; #50; // Sample(116)
        x =              290; #50; // Sample(117)
        x =               47; #50; // Sample(118)
        x =              157; #50; // Sample(119)
        x =              597; #50; // Sample(120)
        x =              314; #50; // Sample(121)
        x =              458; #50; // Sample(122)
        x =              102; #50; // Sample(123)
        x =              -47; #50; // Sample(124)
        x =             -105; #50; // Sample(125)
        x =              338; #50; // Sample(126)
        x =             -133; #50; // Sample(127)
        x =              543; #50; // Sample(128)
        x =              479; #50; // Sample(129)
        x =              307; #50; // Sample(130)
        x =              435; #50; // Sample(131)
        x =              206; #50; // Sample(132)
        x =             -133; #50; // Sample(133)
        x =              174; #50; // Sample(134)
        x =               55; #50; // Sample(135)
        x =              405; #50; // Sample(136)
        x =              216; #50; // Sample(137)
        x =              211; #50; // Sample(138)
        x =               45; #50; // Sample(139)
        x =              -72; #50; // Sample(140)
        x =              131; #50; // Sample(141)
        x =              -23; #50; // Sample(142)
        x =              301; #50; // Sample(143)
        x =              -49; #50; // Sample(144)
        x =             -150; #50; // Sample(145)
        x =              -61; #50; // Sample(146)
        x =              165; #50; // Sample(147)
        x =             -166; #50; // Sample(148)
        x =              -96; #50; // Sample(149)
        x =             -374; #50; // Sample(150)
        x =              -92; #50; // Sample(151)
        x =             -205; #50; // Sample(152)
        x =             -234; #50; // Sample(153)
        x =             -140; #50; // Sample(154)
        x =             -178; #50; // Sample(155)
        x =             -198; #50; // Sample(156)
        x =              354; #50; // Sample(157)
        x =              -29; #50; // Sample(158)
        x =               80; #50; // Sample(159)
        x =               65; #50; // Sample(160)
        x =             -314; #50; // Sample(161)
        x =             -361; #50; // Sample(162)
        x =             -591; #50; // Sample(163)
        x =             -467; #50; // Sample(164)
        x =             -344; #50; // Sample(165)
        x =             -311; #50; // Sample(166)
        x =             -236; #50; // Sample(167)
        x =             -270; #50; // Sample(168)
        x =             -525; #50; // Sample(169)
        x =             -361; #50; // Sample(170)
        x =               30; #50; // Sample(171)
        x =             -351; #50; // Sample(172)
        x =             -464; #50; // Sample(173)
        x =             -332; #50; // Sample(174)
        x =             -214; #50; // Sample(175)
        x =             -342; #50; // Sample(176)
        x =             -341; #50; // Sample(177)
        x =             -314; #50; // Sample(178)
        x =              -13; #50; // Sample(179)
        x =              -67; #50; // Sample(180)
        x =             -354; #50; // Sample(181)
        x =             -339; #50; // Sample(182)
        x =             -512; #50; // Sample(183)
        x =               46; #50; // Sample(184)
        x =             -170; #50; // Sample(185)
        x =             -179; #50; // Sample(186)
        x =              -81; #50; // Sample(187)
        x =             -342; #50; // Sample(188)
        x =             -252; #50; // Sample(189)
        x =              -24; #50; // Sample(190)
        x =             -100; #50; // Sample(191)
        x =             -409; #50; // Sample(192)
        x =             -146; #50; // Sample(193)
        x =               70; #50; // Sample(194)
        x =              242; #50; // Sample(195)
        x =               76; #50; // Sample(196)
        x =              105; #50; // Sample(197)
        x =                5; #50; // Sample(198)
        x =              155; #50; // Sample(199)
        x =              236; #50; // Sample(200)
        x =              -21; #50; // Sample(201)
        x =              366; #50; // Sample(202)
        x =             -132; #50; // Sample(203)
        x =              189; #50; // Sample(204)
        x =              168; #50; // Sample(205)
        x =              538; #50; // Sample(206)
        x =              179; #50; // Sample(207)
        x =              861; #50; // Sample(208)
        x =              208; #50; // Sample(209)
        x =              133; #50; // Sample(210)
        x =              718; #50; // Sample(211)
        x =              280; #50; // Sample(212)
        x =              241; #50; // Sample(213)
        x =              322; #50; // Sample(214)
        x =              107; #50; // Sample(215)
        x =               22; #50; // Sample(216)
        x =              178; #50; // Sample(217)
        x =              312; #50; // Sample(218)
        x =              514; #50; // Sample(219)
        x =              524; #50; // Sample(220)
        x =              381; #50; // Sample(221)
        x =              511; #50; // Sample(222)
        x =              775; #50; // Sample(223)
        x =              393; #50; // Sample(224)
        x =              443; #50; // Sample(225)
        x =              192; #50; // Sample(226)
        x =              466; #50; // Sample(227)
        x =               12; #50; // Sample(228)
        x =              149; #50; // Sample(229)
        x =               35; #50; // Sample(230)
        x =               77; #50; // Sample(231)
        x =              545; #50; // Sample(232)
        x =              111; #50; // Sample(233)
        x =               52; #50; // Sample(234)
        x =              311; #50; // Sample(235)
        x =               36; #50; // Sample(236)
        x =              139; #50; // Sample(237)
        x =              164; #50; // Sample(238)
        x =             -126; #50; // Sample(239)
        x =              -47; #50; // Sample(240)
        x =              365; #50; // Sample(241)
        x =                6; #50; // Sample(242)
        x =              133; #50; // Sample(243)
        x =              184; #50; // Sample(244)
        x =               32; #50; // Sample(245)
        x =              -72; #50; // Sample(246)
        x =              129; #50; // Sample(247)
        x =             -372; #50; // Sample(248)
        x =               80; #50; // Sample(249)
        x =             -567; #50; // Sample(250)
        x =             -423; #50; // Sample(251)
        x =             -279; #50; // Sample(252)
        x =             -228; #50; // Sample(253)
        x =             -536; #50; // Sample(254)
        x =              -90; #50; // Sample(255)
        x =             -264; #50; // Sample(256)
        x =             -469; #50; // Sample(257)
        x =             -496; #50; // Sample(258)
        x =             -460; #50; // Sample(259)
        x =             -443; #50; // Sample(260)
        x =             -314; #50; // Sample(261)
        x =             -304; #50; // Sample(262)
        x =             -408; #50; // Sample(263)
        x =             -315; #50; // Sample(264)
        x =             -423; #50; // Sample(265)
        x =             -265; #50; // Sample(266)
        x =               -2; #50; // Sample(267)
        x =             -130; #50; // Sample(268)
        x =             -368; #50; // Sample(269)
        x =             -256; #50; // Sample(270)
        x =             -307; #50; // Sample(271)
        x =             -350; #50; // Sample(272)
        x =             -320; #50; // Sample(273)
        x =              -38; #50; // Sample(274)
        x =             -342; #50; // Sample(275)
        x =             -190; #50; // Sample(276)
        x =              -95; #50; // Sample(277)
        x =             -395; #50; // Sample(278)
        x =             -470; #50; // Sample(279)
        x =              -21; #50; // Sample(280)
        x =              -77; #50; // Sample(281)
        x =             -235; #50; // Sample(282)
        x =              100; #50; // Sample(283)
        x =              -36; #50; // Sample(284)
        x =             -155; #50; // Sample(285)
        x =             -143; #50; // Sample(286)
        x =             -134; #50; // Sample(287)
        x =             -228; #50; // Sample(288)
        x =              519; #50; // Sample(289)
        x =             -412; #50; // Sample(290)
        x =               91; #50; // Sample(291)
        x =               60; #50; // Sample(292)
        x =             -166; #50; // Sample(293)
        x =               68; #50; // Sample(294)
        x =              189; #50; // Sample(295)
        x =              328; #50; // Sample(296)
        x =              171; #50; // Sample(297)
        x =              278; #50; // Sample(298)
        x =              516; #50; // Sample(299)
        x =              177; #50; // Sample(300)
        x =              103; #50; // Sample(301)
        x =              -46; #50; // Sample(302)
        x =              399; #50; // Sample(303)
        x =              152; #50; // Sample(304)
        x =              530; #50; // Sample(305)
        x =              283; #50; // Sample(306)
        x =              251; #50; // Sample(307)
        x =              177; #50; // Sample(308)
        x =              192; #50; // Sample(309)
        x =               54; #50; // Sample(310)
        x =              411; #50; // Sample(311)
        x =              219; #50; // Sample(312)
        x =              421; #50; // Sample(313)
        x =              -22; #50; // Sample(314)
        x =              362; #50; // Sample(315)
        x =              120; #50; // Sample(316)
        x =               -7; #50; // Sample(317)
        x =              239; #50; // Sample(318)
        x =              394; #50; // Sample(319)
        x =              465; #50; // Sample(320)
        x =              494; #50; // Sample(321)
        x =              177; #50; // Sample(322)
        x =               56; #50; // Sample(323)
        x =              802; #50; // Sample(324)
        x =              108; #50; // Sample(325)
        x =               64; #50; // Sample(326)
        x =              273; #50; // Sample(327)
        x =              -37; #50; // Sample(328)
        x =               24; #50; // Sample(329)
        x =             -156; #50; // Sample(330)
        x =               77; #50; // Sample(331)
        x =             -117; #50; // Sample(332)
        x =              152; #50; // Sample(333)
        x =               95; #50; // Sample(334)
        x =              -97; #50; // Sample(335)
        x =              -53; #50; // Sample(336)
        x =             -108; #50; // Sample(337)
        x =               12; #50; // Sample(338)
        x =             -163; #50; // Sample(339)
        x =               -8; #50; // Sample(340)
        x =             -239; #50; // Sample(341)
        x =               15; #50; // Sample(342)
        x =             -146; #50; // Sample(343)
        x =             -521; #50; // Sample(344)
        x =             -114; #50; // Sample(345)
        x =               12; #50; // Sample(346)
        x =               56; #50; // Sample(347)
        x =             -155; #50; // Sample(348)
        x =               68; #50; // Sample(349)
        x =              -95; #50; // Sample(350)
        x =              160; #50; // Sample(351)
        x =             -199; #50; // Sample(352)
        x =             -169; #50; // Sample(353)
        x =             -187; #50; // Sample(354)
        x =             -172; #50; // Sample(355)
        x =             -127; #50; // Sample(356)
        x =              -89; #50; // Sample(357)
        x =             -480; #50; // Sample(358)
        x =             -542; #50; // Sample(359)
        x =              -47; #50; // Sample(360)
        x =             -117; #50; // Sample(361)
        x =             -459; #50; // Sample(362)
        x =             -306; #50; // Sample(363)
        x =               55; #50; // Sample(364)
        x =             -508; #50; // Sample(365)
        x =             -222; #50; // Sample(366)
        x =             -539; #50; // Sample(367)
        x =             -236; #50; // Sample(368)
        x =             -202; #50; // Sample(369)
        x =             -283; #50; // Sample(370)
        x =              -60; #50; // Sample(371)
        x =             -252; #50; // Sample(372)
        x =               12; #50; // Sample(373)
        x =                9; #50; // Sample(374)
        x =             -235; #50; // Sample(375)
        x =             -118; #50; // Sample(376)
        x =             -110; #50; // Sample(377)
        x =               50; #50; // Sample(378)
        x =              120; #50; // Sample(379)
        x =               54; #50; // Sample(380)
        x =              -73; #50; // Sample(381)
        x =             -227; #50; // Sample(382)
        x =             -282; #50; // Sample(383)
        x =              188; #50; // Sample(384)
        x =              377; #50; // Sample(385)
        x =               71; #50; // Sample(386)
        x =               26; #50; // Sample(387)
        x =              236; #50; // Sample(388)
        x =             -239; #50; // Sample(389)
        x =               47; #50; // Sample(390)
        x =             -262; #50; // Sample(391)
        x =              214; #50; // Sample(392)
        x =              156; #50; // Sample(393)
        x =              229; #50; // Sample(394)
        x =              102; #50; // Sample(395)
        x =             -154; #50; // Sample(396)
        x =              400; #50; // Sample(397)
        x =              103; #50; // Sample(398)
        x =              272; #50; // Sample(399)
        x =              429; #50; // Sample(400)
        x =              368; #50; // Sample(401)
        x =              113; #50; // Sample(402)
        x =              228; #50; // Sample(403)
        x =              243; #50; // Sample(404)
        x =              477; #50; // Sample(405)
        x =              537; #50; // Sample(406)
        x =               97; #50; // Sample(407)
        x =              107; #50; // Sample(408)
        x =              325; #50; // Sample(409)
        x =              299; #50; // Sample(410)
        x =              335; #50; // Sample(411)
        x =               96; #50; // Sample(412)
        x =               37; #50; // Sample(413)
        x =              269; #50; // Sample(414)
        x =              511; #50; // Sample(415)
        x =              389; #50; // Sample(416)
        x =              238; #50; // Sample(417)
        x =              177; #50; // Sample(418)
        x =               26; #50; // Sample(419)
        x =              396; #50; // Sample(420)
        x =              374; #50; // Sample(421)
        x =              167; #50; // Sample(422)
        x =              256; #50; // Sample(423)
        x =              219; #50; // Sample(424)
        x =              325; #50; // Sample(425)
        x =              443; #50; // Sample(426)
        x =             -217; #50; // Sample(427)
        x =               38; #50; // Sample(428)
        x =               63; #50; // Sample(429)
        x =             -182; #50; // Sample(430)
        x =              -16; #50; // Sample(431)
        x =              174; #50; // Sample(432)
        x =             -143; #50; // Sample(433)
        x =             -417; #50; // Sample(434)
        x =             -232; #50; // Sample(435)
        x =               -5; #50; // Sample(436)
        x =             -222; #50; // Sample(437)
        x =               83; #50; // Sample(438)
        x =             -220; #50; // Sample(439)
        x =              -89; #50; // Sample(440)
        x =             -263; #50; // Sample(441)
        x =              -48; #50; // Sample(442)
        x =             -493; #50; // Sample(443)
        x =              112; #50; // Sample(444)
        x =             -253; #50; // Sample(445)
        x =             -252; #50; // Sample(446)
        x =             -507; #50; // Sample(447)
        x =             -249; #50; // Sample(448)
        x =             -273; #50; // Sample(449)
        x =             -497; #50; // Sample(450)
        x =             -164; #50; // Sample(451)
        x =               96; #50; // Sample(452)
        x =              -65; #50; // Sample(453)
        x =             -306; #50; // Sample(454)
        x =             -192; #50; // Sample(455)
        x =             -259; #50; // Sample(456)
        x =             -221; #50; // Sample(457)
        x =             -689; #50; // Sample(458)
        x =             -468; #50; // Sample(459)
        x =             -348; #50; // Sample(460)
        x =             -170; #50; // Sample(461)
        x =             -215; #50; // Sample(462)
        x =             -296; #50; // Sample(463)
        x =             -677; #50; // Sample(464)
        x =             -529; #50; // Sample(465)
        x =                4; #50; // Sample(466)
        x =             -212; #50; // Sample(467)
        x =             -223; #50; // Sample(468)
        x =             -276; #50; // Sample(469)
        x =              351; #50; // Sample(470)
        x =             -312; #50; // Sample(471)
        x =             -194; #50; // Sample(472)
        x =              -49; #50; // Sample(473)
        x =              117; #50; // Sample(474)
        x =             -140; #50; // Sample(475)
        x =               87; #50; // Sample(476)
        x =              110; #50; // Sample(477)
        x =              -10; #50; // Sample(478)
        x =             -287; #50; // Sample(479)
        x =              132; #50; // Sample(480)
        x =               20; #50; // Sample(481)
        x =              313; #50; // Sample(482)
        x =             -119; #50; // Sample(483)
        x =               58; #50; // Sample(484)
        x =              -17; #50; // Sample(485)
        x =             -251; #50; // Sample(486)
        x =              -83; #50; // Sample(487)
        x =             -236; #50; // Sample(488)
        x =              469; #50; // Sample(489)
        x =              213; #50; // Sample(490)
        x =              296; #50; // Sample(491)
        x =              237; #50; // Sample(492)
        x =              423; #50; // Sample(493)
        x =              512; #50; // Sample(494)
        x =              162; #50; // Sample(495)
        x =               67; #50; // Sample(496)
        x =              469; #50; // Sample(497)
        x =              693; #50; // Sample(498)
        x =              236; #50; // Sample(499)
        x =              141; #50; // Sample(500)
        x =                0; #50; // Sample(1)
        x =              183; #50; // Sample(2)
        x =              290; #50; // Sample(3)
        x =              277; #50; // Sample(4)
        x =              150; #50; // Sample(5)
        x =              -39; #50; // Sample(6)
        x =             -212; #50; // Sample(7)
        x =             -297; #50; // Sample(8)
        x =             -260; #50; // Sample(9)
        x =             -115; #50; // Sample(10)
        x =               78; #50; // Sample(11)
        x =              238; #50; // Sample(12)
        x =              300; #50; // Sample(13)
        x =              238; #50; // Sample(14)
        x =               78; #50; // Sample(15)
        x =             -115; #50; // Sample(16)
        x =             -260; #50; // Sample(17)
        x =             -297; #50; // Sample(18)
        x =             -212; #50; // Sample(19)
        x =              -39; #50; // Sample(20)
        x =              150; #50; // Sample(21)
        x =              277; #50; // Sample(22)
        x =              290; #50; // Sample(23)
        x =              183; #50; // Sample(24)
        x =                0; #50; // Sample(25)
        x =             -183; #50; // Sample(26)
        x =             -290; #50; // Sample(27)
        x =             -277; #50; // Sample(28)
        x =             -150; #50; // Sample(29)
        x =               39; #50; // Sample(30)
        x =              212; #50; // Sample(31)
        x =              297; #50; // Sample(32)
        x =              260; #50; // Sample(33)
        x =              115; #50; // Sample(34)
        x =              -78; #50; // Sample(35)
        x =             -238; #50; // Sample(36)
        x =             -300; #50; // Sample(37)
        x =             -238; #50; // Sample(38)
        x =              -78; #50; // Sample(39)
        x =              115; #50; // Sample(40)
        x =              260; #50; // Sample(41)
        x =              297; #50; // Sample(42)
        x =              212; #50; // Sample(43)
        x =               39; #50; // Sample(44)
        x =             -150; #50; // Sample(45)
        x =             -277; #50; // Sample(46)
        x =             -290; #50; // Sample(47)
        x =             -183; #50; // Sample(48)
        x =               -0; #50; // Sample(49)
        x =              183; #50; // Sample(50)
        x =              290; #50; // Sample(51)
        x =              277; #50; // Sample(52)

/*
        x =              150; #50; // Sample(53)
        x =              -39; #50; // Sample(54)
        x =             -212; #50; // Sample(55)
        x =             -297; #50; // Sample(56)
        x =             -260; #50; // Sample(57)
        x =             -115; #50; // Sample(58)
        x =               78; #50; // Sample(59)
        x =              238; #50; // Sample(60)
        x =              300; #50; // Sample(61)
        x =              238; #50; // Sample(62)
        x =               78; #50; // Sample(63)
        x =             -115; #50; // Sample(64)
        x =             -260; #50; // Sample(65)
        x =             -297; #50; // Sample(66)
        x =             -212; #50; // Sample(67)
        x =              -39; #50; // Sample(68)
        x =              150; #50; // Sample(69)
        x =              277; #50; // Sample(70)
        x =              290; #50; // Sample(71)
        x =              183; #50; // Sample(72)
        x =               -0; #50; // Sample(73)
        x =             -183; #50; // Sample(74)
        x =             -290; #50; // Sample(75)
        x =             -277; #50; // Sample(76)
        x =             -150; #50; // Sample(77)
        x =               39; #50; // Sample(78)
        x =              212; #50; // Sample(79)
        x =              297; #50; // Sample(80)
        x =              260; #50; // Sample(81)
        x =              115; #50; // Sample(82)
        x =              -78; #50; // Sample(83)
        x =             -238; #50; // Sample(84)
        x =             -300; #50; // Sample(85)
        x =             -238; #50; // Sample(86)
        x =              -78; #50; // Sample(87)
        x =              115; #50; // Sample(88)
        x =              260; #50; // Sample(89)
        x =              297; #50; // Sample(90)
        x =              212; #50; // Sample(91)
        x =               39; #50; // Sample(92)
        x =             -150; #50; // Sample(93)
        x =             -277; #50; // Sample(94)
        x =             -290; #50; // Sample(95)
        x =             -183; #50; // Sample(96)
        x =               -0; #50; // Sample(97)
        x =              183; #50; // Sample(98)
        x =              290; #50; // Sample(99)
        x =              277; #50; // Sample(100)
        x =              150; #50; // Sample(101)
        x =              -39; #50; // Sample(102)
        x =             -212; #50; // Sample(103)
        x =             -297; #50; // Sample(104)
        x =             -260; #50; // Sample(105)
        x =             -115; #50; // Sample(106)
        x =               78; #50; // Sample(107)
        x =              238; #50; // Sample(108)
        x =              300; #50; // Sample(109)
        x =              238; #50; // Sample(110)
        x =               78; #50; // Sample(111)
        x =             -115; #50; // Sample(112)
        x =             -260; #50; // Sample(113)
        x =             -297; #50; // Sample(114)
        x =             -212; #50; // Sample(115)
        x =              -39; #50; // Sample(116)
        x =              150; #50; // Sample(117)
        x =              277; #50; // Sample(118)
        x =              290; #50; // Sample(119)
        x =              183; #50; // Sample(120)
        x =               -0; #50; // Sample(121)
        x =             -183; #50; // Sample(122)
        x =             -290; #50; // Sample(123)
        x =             -277; #50; // Sample(124)
        x =             -150; #50; // Sample(125)
        x =               39; #50; // Sample(126)
        x =              212; #50; // Sample(127)
        x =              297; #50; // Sample(128)
        x =              260; #50; // Sample(129)
        x =              115; #50; // Sample(130)
        x =              -78; #50; // Sample(131)
        x =             -238; #50; // Sample(132)
        x =             -300; #50; // Sample(133)
        x =             -238; #50; // Sample(134)
        x =              -78; #50; // Sample(135)
        x =              115; #50; // Sample(136)
        x =              260; #50; // Sample(137)
        x =              297; #50; // Sample(138)
        x =              212; #50; // Sample(139)
        x =               39; #50; // Sample(140)
        x =             -150; #50; // Sample(141)
        x =             -277; #50; // Sample(142)
        x =             -290; #50; // Sample(143)
        x =             -183; #50; // Sample(144)
        x =                0; #50; // Sample(145)
        x =              183; #50; // Sample(146)
        x =              290; #50; // Sample(147)
        x =              277; #50; // Sample(148)
        x =              150; #50; // Sample(149)
        x =              -39; #50; // Sample(150)
        x =             -212; #50; // Sample(151)
        x =             -297; #50; // Sample(152)
        x =             -260; #50; // Sample(153)
        x =             -115; #50; // Sample(154)
        x =               78; #50; // Sample(155)
        x =              238; #50; // Sample(156)
        x =              300; #50; // Sample(157)
        x =              238; #50; // Sample(158)
        x =               78; #50; // Sample(159)
        x =             -115; #50; // Sample(160)
        x =             -260; #50; // Sample(161)
        x =             -297; #50; // Sample(162)
        x =             -212; #50; // Sample(163)
        x =              -39; #50; // Sample(164)
        x =              150; #50; // Sample(165)
        x =              277; #50; // Sample(166)
        x =              290; #50; // Sample(167)
        x =              183; #50; // Sample(168)
        x =               -0; #50; // Sample(169)
        x =             -183; #50; // Sample(170)
        x =             -290; #50; // Sample(171)
        x =             -277; #50; // Sample(172)
        x =             -150; #50; // Sample(173)
        x =               39; #50; // Sample(174)
        x =              212; #50; // Sample(175)
        x =              297; #50; // Sample(176)
        x =              260; #50; // Sample(177)
        x =              115; #50; // Sample(178)
        x =              -78; #50; // Sample(179)
        x =             -238; #50; // Sample(180)
        x =             -300; #50; // Sample(181)
        x =             -238; #50; // Sample(182)
        x =              -78; #50; // Sample(183)
        x =              115; #50; // Sample(184)
        x =              260; #50; // Sample(185)
        x =              297; #50; // Sample(186)
        x =              212; #50; // Sample(187)
        x =               39; #50; // Sample(188)
        x =             -150; #50; // Sample(189)
        x =             -277; #50; // Sample(190)
        x =             -290; #50; // Sample(191)
        x =             -183; #50; // Sample(192)
        x =               -0; #50; // Sample(193)
        x =              183; #50; // Sample(194)
        x =              290; #50; // Sample(195)
        x =              277; #50; // Sample(196)
        x =              150; #50; // Sample(197)
        x =              -39; #50; // Sample(198)
        x =             -212; #50; // Sample(199)
        x =             -297; #50; // Sample(200)
        x =             -260; #50; // Sample(201)
        x =             -115; #50; // Sample(202)
        x =               78; #50; // Sample(203)
        x =              238; #50; // Sample(204)
        x =              300; #50; // Sample(205)
        x =              238; #50; // Sample(206)
        x =               78; #50; // Sample(207)
        x =             -115; #50; // Sample(208)
        x =             -260; #50; // Sample(209)
        x =             -297; #50; // Sample(210)
        x =             -212; #50; // Sample(211)
        x =              -39; #50; // Sample(212)
        x =              150; #50; // Sample(213)
        x =              277; #50; // Sample(214)
        x =              290; #50; // Sample(215)
        x =              183; #50; // Sample(216)
        x =                0; #50; // Sample(217)
        x =             -183; #50; // Sample(218)
        x =             -290; #50; // Sample(219)
        x =             -277; #50; // Sample(220)
        x =             -150; #50; // Sample(221)
        x =               39; #50; // Sample(222)
        x =              212; #50; // Sample(223)
        x =              297; #50; // Sample(224)
        x =              260; #50; // Sample(225)
        x =              115; #50; // Sample(226)
        x =              -78; #50; // Sample(227)
        x =             -238; #50; // Sample(228)
        x =             -300; #50; // Sample(229)
        x =             -238; #50; // Sample(230)
        x =              -78; #50; // Sample(231)
        x =              115; #50; // Sample(232)
        x =              260; #50; // Sample(233)
        x =              297; #50; // Sample(234)
        x =              212; #50; // Sample(235)
        x =               39; #50; // Sample(236)
        x =             -150; #50; // Sample(237)
        x =             -277; #50; // Sample(238)
        x =             -290; #50; // Sample(239)
        x =             -183; #50; // Sample(240)
        x =                0; #50; // Sample(241)
        x =              183; #50; // Sample(242)
        x =              290; #50; // Sample(243)
        x =              277; #50; // Sample(244)
        x =              150; #50; // Sample(245)
        x =              -39; #50; // Sample(246)
        x =             -212; #50; // Sample(247)
        x =             -297; #50; // Sample(248)
        x =             -260; #50; // Sample(249)
        x =             -115; #50; // Sample(250)
        x =               78; #50; // Sample(251)
        x =              238; #50; // Sample(252)
        x =              300; #50; // Sample(253)
        x =              238; #50; // Sample(254)
        x =               78; #50; // Sample(255)
        x =             -115; #50; // Sample(256)
        x =             -260; #50; // Sample(257)
        x =             -297; #50; // Sample(258)
        x =             -212; #50; // Sample(259)
        x =              -39; #50; // Sample(260)
        x =              150; #50; // Sample(261)
        x =              277; #50; // Sample(262)
        x =              290; #50; // Sample(263)
        x =              183; #50; // Sample(264)
        x =               -0; #50; // Sample(265)
        x =             -183; #50; // Sample(266)
        x =             -290; #50; // Sample(267)
        x =             -277; #50; // Sample(268)
        x =             -150; #50; // Sample(269)
        x =               39; #50; // Sample(270)
        x =              212; #50; // Sample(271)
        x =              297; #50; // Sample(272)
        x =              260; #50; // Sample(273)
        x =              115; #50; // Sample(274)
        x =              -78; #50; // Sample(275)
        x =             -238; #50; // Sample(276)
        x =             -300; #50; // Sample(277)
        x =             -238; #50; // Sample(278)
        x =              -78; #50; // Sample(279)
        x =              115; #50; // Sample(280)
        x =              260; #50; // Sample(281)
        x =              297; #50; // Sample(282)
        x =              212; #50; // Sample(283)
        x =               39; #50; // Sample(284)
        x =             -150; #50; // Sample(285)
        x =             -277; #50; // Sample(286)
        x =             -290; #50; // Sample(287)
        x =             -183; #50; // Sample(288)
        x =                0; #50; // Sample(289)
        x =              183; #50; // Sample(290)
        x =              290; #50; // Sample(291)
        x =              277; #50; // Sample(292)
        x =              150; #50; // Sample(293)
        x =              -39; #50; // Sample(294)
        x =             -212; #50; // Sample(295)
        x =             -297; #50; // Sample(296)
        x =             -260; #50; // Sample(297)
        x =             -115; #50; // Sample(298)
        x =               78; #50; // Sample(299)
        x =              238; #50; // Sample(300)
        x =              300; #50; // Sample(301)
        x =              238; #50; // Sample(302)
        x =               78; #50; // Sample(303)
        x =             -115; #50; // Sample(304)
        x =             -260; #50; // Sample(305)
        x =             -297; #50; // Sample(306)
        x =             -212; #50; // Sample(307)
        x =              -39; #50; // Sample(308)
        x =              150; #50; // Sample(309)
        x =              277; #50; // Sample(310)
        x =              290; #50; // Sample(311)
        x =              183; #50; // Sample(312)
        x =               -0; #50; // Sample(313)
        x =             -183; #50; // Sample(314)
        x =             -290; #50; // Sample(315)
        x =             -277; #50; // Sample(316)
        x =             -150; #50; // Sample(317)
        x =               39; #50; // Sample(318)
        x =              212; #50; // Sample(319)
        x =              297; #50; // Sample(320)
        x =              260; #50; // Sample(321)
        x =              115; #50; // Sample(322)
        x =              -78; #50; // Sample(323)
        x =             -238; #50; // Sample(324)
        x =             -300; #50; // Sample(325)
        x =             -238; #50; // Sample(326)
        x =              -78; #50; // Sample(327)
        x =              115; #50; // Sample(328)
        x =              260; #50; // Sample(329)
        x =              297; #50; // Sample(330)
        x =              212; #50; // Sample(331)
        x =               39; #50; // Sample(332)
        x =             -150; #50; // Sample(333)
        x =             -277; #50; // Sample(334)
        x =             -290; #50; // Sample(335)
        x =             -183; #50; // Sample(336)
        x =                0; #50; // Sample(337)
        x =              183; #50; // Sample(338)
        x =              290; #50; // Sample(339)
        x =              277; #50; // Sample(340)
        x =              150; #50; // Sample(341)
        x =              -39; #50; // Sample(342)
*/
        $finish;
    end
endmodule
