`timescale 1ns / 1ps

module testbench;

  // All Parameters and Inputs
  // Params
  localparam ORDER = 2;
  localparam FAC = 24;
  localparam BITWIDTH = 32;
  localparam GAINL = 0;
  localparam GAINM = 0;
  localparam HTP = 10;
  // Params End

  reg clk, reset;
  reg signed [BITWIDTH-1:0] x;
  wire signed [BITWIDTH-1:0] y;

  // Instantiate the Unit Under Test (DUT)
  iir_N #(.N(ORDER), .BITWIDTH(BITWIDTH), .FAC(FAC), .GAINL(GAINL), .GAINM(GAINM)) DUT(
    .clk(clk),
    .rst(reset),
    .x(x),
    .y(y)
  );

  // Generate clock with 2*htp period
  initial clk = 0;
  always #HTP clk = ~clk;
  
  always @(posedge(clk)) $display("x = %.0f, y = %.0f", x, y);

  initial begin
    // Begin Init Sequence
    x = {(BITWIDTH-1){1'b0}};
    reset = 1;
    clk = 0;
    clk = 1;
    #10;
    reset = 0;
    #20;

    // Input Stimuli - Python Script adds input lines using Stimuli and Stimuli End comment
//{
    // Stimuli
		#(2*HTP); x = 25;
		#(2*HTP); x = 10;
		#(2*HTP); x = 25;
		#(2*HTP); x = 10;
		#(2*HTP); x = 67;
		#(2*HTP); x = -56;
		#(2*HTP); x = 19;
		#(2*HTP); x = 28;
		#(2*HTP); x = 160;
		#(2*HTP); x = 39;
		#(2*HTP); x = 142;
		#(2*HTP); x = 151;
		#(2*HTP); x = 117;
		#(2*HTP); x = 294;
		#(2*HTP); x = 199;
		#(2*HTP); x = 363;
		#(2*HTP); x = 100;
		#(2*HTP); x = 525;
		#(2*HTP); x = 78;
		#(2*HTP); x = 195;
		#(2*HTP); x = -19;
		#(2*HTP); x = 147;
		#(2*HTP); x = 515;
		#(2*HTP); x = 373;
		#(2*HTP); x = 110;
		#(2*HTP); x = 389;
		#(2*HTP); x = 161;
		#(2*HTP); x = -98;
		#(2*HTP); x = 198;
		#(2*HTP); x = 673;
		#(2*HTP); x = 338;
		#(2*HTP); x = -79;
		#(2*HTP); x = 424;
		#(2*HTP); x = 653;
		#(2*HTP); x = 269;
		#(2*HTP); x = 241;
		#(2*HTP); x = 374;
		#(2*HTP); x = 92;
		#(2*HTP); x = 296;
		#(2*HTP); x = 707;
		#(2*HTP); x = 46;
		#(2*HTP); x = 212;
		#(2*HTP); x = 262;
		#(2*HTP); x = 251;
		#(2*HTP); x = 315;
		#(2*HTP); x = 94;
		#(2*HTP); x = -26;
		#(2*HTP); x = 84;
		#(2*HTP); x = -286;
		#(2*HTP); x = 18;
		#(2*HTP); x = 459;
		#(2*HTP); x = -86;
		#(2*HTP); x = 70;
		#(2*HTP); x = 77;
		#(2*HTP); x = 38;
		#(2*HTP); x = -44;
		#(2*HTP); x = -200;
		#(2*HTP); x = -27;
		#(2*HTP); x = -67;
		#(2*HTP); x = -100;
		#(2*HTP); x = -33;
		#(2*HTP); x = -199;
		#(2*HTP); x = -407;
		#(2*HTP); x = -343;
		#(2*HTP); x = -78;
		#(2*HTP); x = -28;
		#(2*HTP); x = -358;
		#(2*HTP); x = -503;
		#(2*HTP); x = -454;
		#(2*HTP); x = -75;
		#(2*HTP); x = -101;
		#(2*HTP); x = -133;
		#(2*HTP); x = -103;
		#(2*HTP); x = -299;
		#(2*HTP); x = -267;
		#(2*HTP); x = -161;
		#(2*HTP); x = -123;
		#(2*HTP); x = 191;
		#(2*HTP); x = -482;
		#(2*HTP); x = -272;
		#(2*HTP); x = -206;
		#(2*HTP); x = -506;
		#(2*HTP); x = -562;
		#(2*HTP); x = -238;
		#(2*HTP); x = -396;
		#(2*HTP); x = -249;
		#(2*HTP); x = -421;
		#(2*HTP); x = -245;
		#(2*HTP); x = -193;
		#(2*HTP); x = -624;
		#(2*HTP); x = -37;
		#(2*HTP); x = -554;
		#(2*HTP); x = -101;
		#(2*HTP); x = -129;
		#(2*HTP); x = -70;
		#(2*HTP); x = 197;
		#(2*HTP); x = -374;
		#(2*HTP); x = -191;
		#(2*HTP); x = -186;
		#(2*HTP); x = 278;
		#(2*HTP); x = 253;
		#(2*HTP); x = 156;
		#(2*HTP); x = -260;
		#(2*HTP); x = -30;
		#(2*HTP); x = 179;
		#(2*HTP); x = 164;
		#(2*HTP); x = -10;
		#(2*HTP); x = 423;
		#(2*HTP); x = 39;
		#(2*HTP); x = 241;
		#(2*HTP); x = 568;
		#(2*HTP); x = 532;
		#(2*HTP); x = 174;
		#(2*HTP); x = 371;
		#(2*HTP); x = 562;
		#(2*HTP); x = 66;
		#(2*HTP); x = 445;
		#(2*HTP); x = 628;
		#(2*HTP); x = 471;
		#(2*HTP); x = 522;
		#(2*HTP); x = 290;
		#(2*HTP); x = 47;
		#(2*HTP); x = 157;
		#(2*HTP); x = 597;
		#(2*HTP); x = 314;
		#(2*HTP); x = 458;
		#(2*HTP); x = 102;
		#(2*HTP); x = -47;
		#(2*HTP); x = -105;
		#(2*HTP); x = 338;
		#(2*HTP); x = -133;
		#(2*HTP); x = 543;
		#(2*HTP); x = 479;
		#(2*HTP); x = 307;
		#(2*HTP); x = 435;
		#(2*HTP); x = 206;
		#(2*HTP); x = -133;
		#(2*HTP); x = 174;
		#(2*HTP); x = 55;
		#(2*HTP); x = 405;
		#(2*HTP); x = 216;
		#(2*HTP); x = 211;
		#(2*HTP); x = 45;
		#(2*HTP); x = -72;
		#(2*HTP); x = 131;
		#(2*HTP); x = -23;
		#(2*HTP); x = 301;
		#(2*HTP); x = -49;
		#(2*HTP); x = -150;
		#(2*HTP); x = -61;
		#(2*HTP); x = 165;
		#(2*HTP); x = -166;
		#(2*HTP); x = -96;
		#(2*HTP); x = -374;
		#(2*HTP); x = -92;
		#(2*HTP); x = -205;
		#(2*HTP); x = -234;
		#(2*HTP); x = -140;
		#(2*HTP); x = -178;
		#(2*HTP); x = -198;
		#(2*HTP); x = 354;
		#(2*HTP); x = -29;
		#(2*HTP); x = 80;
		#(2*HTP); x = 65;
		#(2*HTP); x = -314;
		#(2*HTP); x = -361;
		#(2*HTP); x = -591;
		#(2*HTP); x = -467;
		#(2*HTP); x = -344;
		#(2*HTP); x = -311;
		#(2*HTP); x = -236;
		#(2*HTP); x = -270;
		#(2*HTP); x = -525;
		#(2*HTP); x = -361;
		#(2*HTP); x = 30;
		#(2*HTP); x = -351;
		#(2*HTP); x = -464;
		#(2*HTP); x = -332;
		#(2*HTP); x = -214;
		#(2*HTP); x = -342;
		#(2*HTP); x = -341;
		#(2*HTP); x = -314;
		#(2*HTP); x = -13;
		#(2*HTP); x = -67;
		#(2*HTP); x = -354;
		#(2*HTP); x = -339;
		#(2*HTP); x = -512;
		#(2*HTP); x = 46;
		#(2*HTP); x = -170;
		#(2*HTP); x = -179;
		#(2*HTP); x = -81;
		#(2*HTP); x = -342;
		#(2*HTP); x = -252;
		#(2*HTP); x = -24;
		#(2*HTP); x = -100;
		#(2*HTP); x = -409;
		#(2*HTP); x = -146;
		#(2*HTP); x = 70;
		#(2*HTP); x = 242;
		#(2*HTP); x = 76;
		#(2*HTP); x = 105;
		#(2*HTP); x = 5;
		#(2*HTP); x = 155;
		#(2*HTP); x = 236;
		#(2*HTP); x = -21;
		#(2*HTP); x = 366;
		#(2*HTP); x = -132;
		#(2*HTP); x = 189;
		#(2*HTP); x = 168;
		#(2*HTP); x = 538;
		#(2*HTP); x = 179;
		#(2*HTP); x = 861;
		#(2*HTP); x = 208;
		#(2*HTP); x = 133;
		#(2*HTP); x = 718;
		#(2*HTP); x = 280;
		#(2*HTP); x = 241;
		#(2*HTP); x = 322;
		#(2*HTP); x = 107;
		#(2*HTP); x = 22;
		#(2*HTP); x = 178;
		#(2*HTP); x = 312;
		#(2*HTP); x = 514;
		#(2*HTP); x = 524;
		#(2*HTP); x = 381;
		#(2*HTP); x = 511;
		#(2*HTP); x = 775;
		#(2*HTP); x = 393;
		#(2*HTP); x = 443;
		#(2*HTP); x = 192;
		#(2*HTP); x = 466;
		#(2*HTP); x = 12;
		#(2*HTP); x = 149;
		#(2*HTP); x = 35;
		#(2*HTP); x = 77;
		#(2*HTP); x = 545;
		#(2*HTP); x = 111;
		#(2*HTP); x = 52;
		#(2*HTP); x = 311;
		#(2*HTP); x = 36;
		#(2*HTP); x = 139;
		#(2*HTP); x = 164;
		#(2*HTP); x = -126;
		#(2*HTP); x = -47;
		#(2*HTP); x = 365;
		#(2*HTP); x = 6;
		#(2*HTP); x = 133;
		#(2*HTP); x = 184;
		#(2*HTP); x = 32;
		#(2*HTP); x = -72;
		#(2*HTP); x = 129;
		#(2*HTP); x = -372;
		#(2*HTP); x = 80;
		#(2*HTP); x = -567;
		#(2*HTP); x = -423;
		#(2*HTP); x = -279;
		#(2*HTP); x = -228;
		#(2*HTP); x = -536;
		#(2*HTP); x = -90;
		#(2*HTP); x = -264;
		#(2*HTP); x = -469;
		#(2*HTP); x = -496;
		#(2*HTP); x = -460;
		#(2*HTP); x = -443;
		#(2*HTP); x = -314;
		#(2*HTP); x = -304;
		#(2*HTP); x = -408;
		#(2*HTP); x = -315;
		#(2*HTP); x = -423;
		#(2*HTP); x = -265;
		#(2*HTP); x = -2;
		#(2*HTP); x = -130;
		#(2*HTP); x = -368;
		#(2*HTP); x = -256;
		#(2*HTP); x = -307;
		#(2*HTP); x = -350;
		#(2*HTP); x = -320;
		#(2*HTP); x = -38;
		#(2*HTP); x = -342;
		#(2*HTP); x = -190;
		#(2*HTP); x = -95;
		#(2*HTP); x = -395;
		#(2*HTP); x = -470;
		#(2*HTP); x = -21;
		#(2*HTP); x = -77;
		#(2*HTP); x = -235;
		#(2*HTP); x = 100;
		#(2*HTP); x = -36;
		#(2*HTP); x = -155;
		#(2*HTP); x = -143;
		#(2*HTP); x = -134;
		#(2*HTP); x = -228;
		#(2*HTP); x = 519;
		#(2*HTP); x = -412;
		#(2*HTP); x = 91;
		#(2*HTP); x = 60;
		#(2*HTP); x = -166;
		#(2*HTP); x = 68;
		#(2*HTP); x = 189;
		#(2*HTP); x = 328;
		#(2*HTP); x = 171;
		#(2*HTP); x = 278;
		#(2*HTP); x = 516;
		#(2*HTP); x = 177;
		#(2*HTP); x = 103;
		#(2*HTP); x = -46;
		#(2*HTP); x = 399;
		#(2*HTP); x = 152;
		#(2*HTP); x = 530;
		#(2*HTP); x = 283;
		#(2*HTP); x = 251;
		#(2*HTP); x = 177;
		#(2*HTP); x = 192;
		#(2*HTP); x = 54;
		#(2*HTP); x = 411;
		#(2*HTP); x = 219;
		#(2*HTP); x = 421;
		#(2*HTP); x = -22;
		#(2*HTP); x = 362;
		#(2*HTP); x = 120;
		#(2*HTP); x = -7;
		#(2*HTP); x = 239;
		#(2*HTP); x = 394;
		#(2*HTP); x = 465;
		#(2*HTP); x = 494;
		#(2*HTP); x = 177;
		#(2*HTP); x = 56;
		#(2*HTP); x = 802;
		#(2*HTP); x = 108;
		#(2*HTP); x = 64;
		#(2*HTP); x = 273;
		#(2*HTP); x = -37;
		#(2*HTP); x = 24;
		#(2*HTP); x = -156;
		#(2*HTP); x = 77;
		#(2*HTP); x = -117;
		#(2*HTP); x = 152;
		#(2*HTP); x = 95;
		#(2*HTP); x = -97;
		#(2*HTP); x = -53;
		#(2*HTP); x = -108;
		#(2*HTP); x = 12;
		#(2*HTP); x = -163;
		#(2*HTP); x = -8;
		#(2*HTP); x = -239;
		#(2*HTP); x = 15;
		#(2*HTP); x = -146;
		#(2*HTP); x = -521;
		#(2*HTP); x = -114;
		#(2*HTP); x = 12;
		#(2*HTP); x = 56;
		#(2*HTP); x = -155;
		#(2*HTP); x = 68;
		#(2*HTP); x = -95;
		#(2*HTP); x = 160;
		#(2*HTP); x = -199;
		#(2*HTP); x = -169;
		#(2*HTP); x = -187;
		#(2*HTP); x = -172;
		#(2*HTP); x = -127;
		#(2*HTP); x = -89;
		#(2*HTP); x = -480;
		#(2*HTP); x = -542;
		#(2*HTP); x = -47;
		#(2*HTP); x = -117;
		#(2*HTP); x = -459;
		#(2*HTP); x = -306;
		#(2*HTP); x = 55;
		#(2*HTP); x = -508;
		#(2*HTP); x = -222;
		#(2*HTP); x = -539;
		#(2*HTP); x = -236;
		#(2*HTP); x = -202;
		#(2*HTP); x = -283;
		#(2*HTP); x = -60;
		#(2*HTP); x = -252;
		#(2*HTP); x = 12;
		#(2*HTP); x = 9;
		#(2*HTP); x = -235;
		#(2*HTP); x = -118;
		#(2*HTP); x = -110;
		#(2*HTP); x = 50;
		#(2*HTP); x = 120;
		#(2*HTP); x = 54;
		#(2*HTP); x = -73;
		#(2*HTP); x = -227;
		#(2*HTP); x = -282;
		#(2*HTP); x = 188;
		#(2*HTP); x = 377;
		#(2*HTP); x = 71;
		#(2*HTP); x = 26;
		#(2*HTP); x = 236;
		#(2*HTP); x = -239;
		#(2*HTP); x = 47;
		#(2*HTP); x = -262;
		#(2*HTP); x = 214;
		#(2*HTP); x = 156;
		#(2*HTP); x = 229;
		#(2*HTP); x = 102;
		#(2*HTP); x = -154;
		#(2*HTP); x = 400;
		#(2*HTP); x = 103;
		#(2*HTP); x = 272;
		#(2*HTP); x = 429;
		#(2*HTP); x = 368;
		#(2*HTP); x = 113;
		#(2*HTP); x = 228;
		#(2*HTP); x = 243;
		#(2*HTP); x = 477;
		#(2*HTP); x = 537;
		#(2*HTP); x = 97;
		#(2*HTP); x = 107;
		#(2*HTP); x = 325;
		#(2*HTP); x = 299;
		#(2*HTP); x = 335;
		#(2*HTP); x = 96;
		#(2*HTP); x = 37;
		#(2*HTP); x = 269;
		#(2*HTP); x = 511;
		#(2*HTP); x = 389;
		#(2*HTP); x = 238;
		#(2*HTP); x = 177;
		#(2*HTP); x = 26;
		#(2*HTP); x = 396;
		#(2*HTP); x = 374;
		#(2*HTP); x = 167;
		#(2*HTP); x = 256;
		#(2*HTP); x = 219;
		#(2*HTP); x = 325;
		#(2*HTP); x = 443;
		#(2*HTP); x = -217;
		#(2*HTP); x = 38;
		#(2*HTP); x = 63;
		#(2*HTP); x = -182;
		#(2*HTP); x = -16;
		#(2*HTP); x = 174;
		#(2*HTP); x = -143;
		#(2*HTP); x = -417;
		#(2*HTP); x = -232;
		#(2*HTP); x = -5;
		#(2*HTP); x = -222;
		#(2*HTP); x = 83;
		#(2*HTP); x = -220;
		#(2*HTP); x = -89;
		#(2*HTP); x = -263;
		#(2*HTP); x = -48;
		#(2*HTP); x = -493;
		#(2*HTP); x = 112;
		#(2*HTP); x = -253;
		#(2*HTP); x = -252;
		#(2*HTP); x = -507;
		#(2*HTP); x = -249;
		#(2*HTP); x = -273;
		#(2*HTP); x = -497;
		#(2*HTP); x = -164;
		#(2*HTP); x = 96;
		#(2*HTP); x = -65;
		#(2*HTP); x = -306;
		#(2*HTP); x = -192;
		#(2*HTP); x = -259;
		#(2*HTP); x = -221;
		#(2*HTP); x = -689;
		#(2*HTP); x = -468;
		#(2*HTP); x = -348;
		#(2*HTP); x = -170;
		#(2*HTP); x = -215;
		#(2*HTP); x = -296;
		#(2*HTP); x = -677;
		#(2*HTP); x = -529;
		#(2*HTP); x = 4;
		#(2*HTP); x = -212;
		#(2*HTP); x = -223;
		#(2*HTP); x = -276;
		#(2*HTP); x = 351;
		#(2*HTP); x = -312;
		#(2*HTP); x = -194;
		#(2*HTP); x = -49;
		#(2*HTP); x = 117;
		#(2*HTP); x = -140;
		#(2*HTP); x = 87;
		#(2*HTP); x = 110;
		#(2*HTP); x = -10;
		#(2*HTP); x = -287;
		#(2*HTP); x = 132;
		#(2*HTP); x = 20;
		#(2*HTP); x = 313;
		#(2*HTP); x = -119;
		#(2*HTP); x = 58;
		#(2*HTP); x = -17;
		#(2*HTP); x = -251;
		#(2*HTP); x = -83;
		#(2*HTP); x = -236;
		#(2*HTP); x = 469;
		#(2*HTP); x = 213;
		#(2*HTP); x = 296;
		#(2*HTP); x = 237;
		#(2*HTP); x = 423;
		#(2*HTP); x = 512;
		#(2*HTP); x = 162;
		#(2*HTP); x = 67;
		#(2*HTP); x = 469;
		#(2*HTP); x = 693;
		#(2*HTP); x = 236;
		#(2*HTP); x = 141;
		#(2*HTP); x = 0;
		#(2*HTP); x = 183;
		#(2*HTP); x = 290;
		#(2*HTP); x = 277;
		#(2*HTP); x = 150;
		#(2*HTP); x = -39;
		#(2*HTP); x = -212;
		#(2*HTP); x = -297;
		#(2*HTP); x = -260;
		#(2*HTP); x = -115;
		#(2*HTP); x = 78;
		#(2*HTP); x = 238;
		#(2*HTP); x = 300;
		#(2*HTP); x = 238;
		#(2*HTP); x = 78;
		#(2*HTP); x = -115;
		#(2*HTP); x = -260;
		#(2*HTP); x = -297;
		#(2*HTP); x = -212;
		#(2*HTP); x = -39;
		#(2*HTP); x = 150;
		#(2*HTP); x = 277;
		#(2*HTP); x = 290;
		#(2*HTP); x = 183;
		#(2*HTP); x = 0;
		#(2*HTP); x = -183;
		#(2*HTP); x = -290;
		#(2*HTP); x = -277;
		#(2*HTP); x = -150;
		#(2*HTP); x = 39;
		#(2*HTP); x = 212;
		#(2*HTP); x = 297;
		#(2*HTP); x = 260;
		#(2*HTP); x = 115;
		#(2*HTP); x = -78;
		#(2*HTP); x = -238;
		#(2*HTP); x = -300;
		#(2*HTP); x = -238;
		#(2*HTP); x = -78;
		#(2*HTP); x = 115;
		#(2*HTP); x = 260;
		#(2*HTP); x = 297;
		#(2*HTP); x = 212;
		#(2*HTP); x = 39;
		#(2*HTP); x = -150;
		#(2*HTP); x = -277;
		#(2*HTP); x = -290;
		#(2*HTP); x = -183;
		#(2*HTP); x = 0;
		#(2*HTP); x = 183;
		#(2*HTP); x = 290;
		#(2*HTP); x = 277;
    // Stimuli End
//}
    $finish;
  end
endmodule